module SA32(clk, rstn, activation, weight, control,c_out0,c_out1,c_out2,c_out3,c_out4,c_out5,c_out6,c_out7,c_out8,c_out9,c_out10,c_out11,c_out12,c_out13,c_out14,c_out15,c_out16,c_out17,c_out18,c_out19,c_out20,c_out21,c_out22,c_out23,c_out24,c_out25,c_out26,c_out27,c_out28,c_out29,c_out30,c_out31,out_act,out_weight);
parameter WIDTH = 8;
parameter C_WIDTH = 32;

input clk,rstn;
input [32*WIDTH-1:0] activation;
input [32*WIDTH-1:0] weight;
input control;
output [32*C_WIDTH-1:0] c_out0;
output [32*C_WIDTH-1:0] c_out1;
output [32*C_WIDTH-1:0] c_out2;
output [32*C_WIDTH-1:0] c_out3;
output [32*C_WIDTH-1:0] c_out4;
output [32*C_WIDTH-1:0] c_out5;
output [32*C_WIDTH-1:0] c_out6;
output [32*C_WIDTH-1:0] c_out7;
output [32*C_WIDTH-1:0] c_out8;
output [32*C_WIDTH-1:0] c_out9;
output [32*C_WIDTH-1:0] c_out10;
output [32*C_WIDTH-1:0] c_out11;
output [32*C_WIDTH-1:0] c_out12;
output [32*C_WIDTH-1:0] c_out13;
output [32*C_WIDTH-1:0] c_out14;
output [32*C_WIDTH-1:0] c_out15;
output [32*C_WIDTH-1:0] c_out16;
output [32*C_WIDTH-1:0] c_out17;
output [32*C_WIDTH-1:0] c_out18;
output [32*C_WIDTH-1:0] c_out19;
output [32*C_WIDTH-1:0] c_out20;
output [32*C_WIDTH-1:0] c_out21;
output [32*C_WIDTH-1:0] c_out22;
output [32*C_WIDTH-1:0] c_out23;
output [32*C_WIDTH-1:0] c_out24;
output [32*C_WIDTH-1:0] c_out25;
output [32*C_WIDTH-1:0] c_out26;
output [32*C_WIDTH-1:0] c_out27;
output [32*C_WIDTH-1:0] c_out28;
output [32*C_WIDTH-1:0] c_out29;
output [32*C_WIDTH-1:0] c_out30;
output [32*C_WIDTH-1:0] c_out31;
output [32*WIDTH-1:0] out_act;
output [32*WIDTH-1:0] out_weight;


wire [16*WIDTH-1:0] act_0;
wire [16*WIDTH-1:0] act_1;
wire [16*WIDTH-1:0] weight_0;
wire [16*WIDTH-1:0] weight_1;

wire [16*WIDTH-1:0] outact_0;
wire [16*WIDTH-1:0] outact_1;
wire [16*WIDTH-1:0] outweight_0;
wire [16*WIDTH-1:0] outweight_1;

wire [16*WIDTH-1:0] act0_1;
wire [16*WIDTH-1:0] act2_3;
wire [16*WIDTH-1:0] weight0_2;
wire [16*WIDTH-1:0] weight1_3;
wire [32*C_WIDTH-1:0] out_0;
wire [32*C_WIDTH-1:0] out_1;
wire [32*C_WIDTH-1:0] out_2;
wire [32*C_WIDTH-1:0] out_3;
wire [32*C_WIDTH-1:0] out_4;
wire [32*C_WIDTH-1:0] out_5;
wire [32*C_WIDTH-1:0] out_6;
wire [32*C_WIDTH-1:0] out_7;
wire [32*C_WIDTH-1:0] out_8;
wire [32*C_WIDTH-1:0] out_9;
wire [32*C_WIDTH-1:0] out_10;
wire [32*C_WIDTH-1:0] out_11;
wire [32*C_WIDTH-1:0] out_12;
wire [32*C_WIDTH-1:0] out_13;
wire [32*C_WIDTH-1:0] out_14;
wire [32*C_WIDTH-1:0] out_15;
wire [32*C_WIDTH-1:0] out_16;
wire [32*C_WIDTH-1:0] out_17;
wire [32*C_WIDTH-1:0] out_18;
wire [32*C_WIDTH-1:0] out_19;
wire [32*C_WIDTH-1:0] out_20;
wire [32*C_WIDTH-1:0] out_21;
wire [32*C_WIDTH-1:0] out_22;
wire [32*C_WIDTH-1:0] out_23;
wire [32*C_WIDTH-1:0] out_24;
wire [32*C_WIDTH-1:0] out_25;
wire [32*C_WIDTH-1:0] out_26;
wire [32*C_WIDTH-1:0] out_27;
wire [32*C_WIDTH-1:0] out_28;
wire [32*C_WIDTH-1:0] out_29;
wire [32*C_WIDTH-1:0] out_30;
wire [32*C_WIDTH-1:0] out_31;

assign {act_0,act_1} = activation;
assign {weight_0,weight_1} = weight;

SA16 SA16_0 (.clk(clk),.rstn(rstn),.activation(act_0),.weight(weight_0),.out_act(act0_1),.out_weight(weight0_2),.control(control),.c_out0(out_0),.c_out1(out_1),.c_out2(out_2),.c_out3(out_3),.c_out4(out_4),.c_out5(out_5),.c_out6(out_6),.c_out7(out_7));
SA16 SA16_1 (.clk(clk),.rstn(rstn),.activation(act0_1),.weight(weight_1),.out_act(outact_0),.out_weight(weight1_3),.control(control),.c_out0(out_8),.c_out1(out_9),.c_out2(out_10),.c_out3(out_11),.c_out4(out_12),.c_out5(out_13),.c_out6(out_14),.c_out7(out_15));
SA16 SA16_2 (.clk(clk),.rstn(rstn),.activation(act_1),.weight(weight0_2),.out_act(act2_3),.out_weight(outweight_0),.control(control),.c_out0(out_16),.c_out1(out_17),.c_out2(out_18),.c_out3(out_19),.c_out4(out_20),.c_out5(out_21),.c_out6(out_22),.c_out7(out_23));
SA16 SA16_3 (.clk(clk),.rstn(rstn),.activation(act2_3),.weight(weight1_3),.out_act(outact_1),.out_weight(outweight_1),.control(control),.c_out0(out_24),.c_out1(out_25),.c_out2(out_26),.c_out3(out_27),.c_out4(out_28),.c_out5(out_29),.c_out6(out_30),.c_out7(out_31));

assign out_act = {outact_0,outact_1};
assign out_weight = {outweight_0,outweight_1};

assign c_out0 = out_0;
assign c_out1 = out_1;
assign c_out2 = out_2;
assign c_out3 = out_3;
assign c_out4 = out_4;
assign c_out5 = out_5;
assign c_out6 = out_6;
assign c_out7 = out_7;
assign c_out8 = out_8;
assign c_out9 = out_9;
assign c_out10 = out_10;
assign c_out11 = out_11;
assign c_out12 = out_12;
assign c_out13 = out_13;
assign c_out14 = out_14;
assign c_out15 = out_15;
assign c_out16 = out_16;
assign c_out17 = out_17;
assign c_out18 = out_18;
assign c_out19 = out_19;
assign c_out20 = out_20;
assign c_out21 = out_21;
assign c_out22 = out_22;
assign c_out23 = out_23;
assign c_out24 = out_24;
assign c_out25 = out_25;
assign c_out26 = out_26;
assign c_out27 = out_27;
assign c_out28 = out_28;
assign c_out29 = out_29;
assign c_out30 = out_30;
assign c_out31 = out_31;

endmodule
