module SA256(clk, rstn, activation, weight, control ,c_out0,c_out1,c_out2,c_out3,c_out4,c_out5,c_out6,c_out7,c_out8,c_out9,c_out10,c_out11,c_out12,c_out13,c_out14,c_out15,c_out16,c_out17,c_out18,c_out19,c_out20,c_out21,c_out22,c_out23,c_out24,c_out25,c_out26,c_out27,c_out28,c_out29,c_out30,c_out31,c_out32,c_out33,c_out34,c_out35,c_out36,c_out37,c_out38,c_out39,c_out40,c_out41,c_out42,c_out43,c_out44,c_out45,c_out46,c_out47,c_out48,c_out49,c_out50,c_out51,c_out52,c_out53,c_out54,c_out55,c_out56,c_out57,c_out58,c_out59,c_out60,c_out61,c_out62,c_out63,c_out64,c_out65,c_out66,c_out67,c_out68,c_out69,c_out70,c_out71,c_out72,c_out73,c_out74,c_out75,c_out76,c_out77,c_out78,c_out79,c_out80,c_out81,c_out82,c_out83,c_out84,c_out85,c_out86,c_out87,c_out88,c_out89,c_out90,c_out91,c_out92,c_out93,c_out94,c_out95,c_out96,c_out97,c_out98,c_out99,c_out100,c_out101,c_out102,c_out103,c_out104,c_out105,c_out106,c_out107,c_out108,c_out109,c_out110,c_out111,c_out112,c_out113,c_out114,c_out115,c_out116,c_out117,c_out118,c_out119,c_out120,c_out121,c_out122,c_out123,c_out124,c_out125,c_out126,c_out127,c_out128,c_out129,c_out130,c_out131,c_out132,c_out133,c_out134,c_out135,c_out136,c_out137,c_out138,c_out139,c_out140,c_out141,c_out142,c_out143,c_out144,c_out145,c_out146,c_out147,c_out148,c_out149,c_out150,c_out151,c_out152,c_out153,c_out154,c_out155,c_out156,c_out157,c_out158,c_out159,c_out160,c_out161,c_out162,c_out163,c_out164,c_out165,c_out166,c_out167,c_out168,c_out169,c_out170,c_out171,c_out172,c_out173,c_out174,c_out175,c_out176,c_out177,c_out178,c_out179,c_out180,c_out181,c_out182,c_out183,c_out184,c_out185,c_out186,c_out187,c_out188,c_out189,c_out190,c_out191,c_out192,c_out193,c_out194,c_out195,c_out196,c_out197,c_out198,c_out199,c_out200,c_out201,c_out202,c_out203,c_out204,c_out205,c_out206,c_out207,c_out208,c_out209,c_out210,c_out211,c_out212,c_out213,c_out214,c_out215,c_out216,c_out217,c_out218,c_out219,c_out220,c_out221,c_out222,c_out223,c_out224,c_out225,c_out226,c_out227,c_out228,c_out229,c_out230,c_out231,c_out232,c_out233,c_out234,c_out235,c_out236,c_out237,c_out238,c_out239,c_out240,c_out241,c_out242,c_out243,c_out244,c_out245,c_out246,c_out247,c_out248,c_out249,c_out250,c_out251,c_out252,c_out253,c_out254,c_out255,c_out256,c_out257,c_out258,c_out259,c_out260,c_out261,c_out262,c_out263,c_out264,c_out265,c_out266,c_out267,c_out268,c_out269,c_out270,c_out271,c_out272,c_out273,c_out274,c_out275,c_out276,c_out277,c_out278,c_out279,c_out280,c_out281,c_out282,c_out283,c_out284,c_out285,c_out286,c_out287,c_out288,c_out289,c_out290,c_out291,c_out292,c_out293,c_out294,c_out295,c_out296,c_out297,c_out298,c_out299,c_out300,c_out301,c_out302,c_out303,c_out304,c_out305,c_out306,c_out307,c_out308,c_out309,c_out310,c_out311,c_out312,c_out313,c_out314,c_out315,c_out316,c_out317,c_out318,c_out319,c_out320,c_out321,c_out322,c_out323,c_out324,c_out325,c_out326,c_out327,c_out328,c_out329,c_out330,c_out331,c_out332,c_out333,c_out334,c_out335,c_out336,c_out337,c_out338,c_out339,c_out340,c_out341,c_out342,c_out343,c_out344,c_out345,c_out346,c_out347,c_out348,c_out349,c_out350,c_out351,c_out352,c_out353,c_out354,c_out355,c_out356,c_out357,c_out358,c_out359,c_out360,c_out361,c_out362,c_out363,c_out364,c_out365,c_out366,c_out367,c_out368,c_out369,c_out370,c_out371,c_out372,c_out373,c_out374,c_out375,c_out376,c_out377,c_out378,c_out379,c_out380,c_out381,c_out382,c_out383,c_out384,c_out385,c_out386,c_out387,c_out388,c_out389,c_out390,c_out391,c_out392,c_out393,c_out394,c_out395,c_out396,c_out397,c_out398,c_out399,c_out400,c_out401,c_out402,c_out403,c_out404,c_out405,c_out406,c_out407,c_out408,c_out409,c_out410,c_out411,c_out412,c_out413,c_out414,c_out415,c_out416,c_out417,c_out418,c_out419,c_out420,c_out421,c_out422,c_out423,c_out424,c_out425,c_out426,c_out427,c_out428,c_out429,c_out430,c_out431,c_out432,c_out433,c_out434,c_out435,c_out436,c_out437,c_out438,c_out439,c_out440,c_out441,c_out442,c_out443,c_out444,c_out445,c_out446,c_out447,c_out448,c_out449,c_out450,c_out451,c_out452,c_out453,c_out454,c_out455,c_out456,c_out457,c_out458,c_out459,c_out460,c_out461,c_out462,c_out463,c_out464,c_out465,c_out466,c_out467,c_out468,c_out469,c_out470,c_out471,c_out472,c_out473,c_out474,c_out475,c_out476,c_out477,c_out478,c_out479,c_out480,c_out481,c_out482,c_out483,c_out484,c_out485,c_out486,c_out487,c_out488,c_out489,c_out490,c_out491,c_out492,c_out493,c_out494,c_out495,c_out496,c_out497,c_out498,c_out499,c_out500,c_out501,c_out502,c_out503,c_out504,c_out505,c_out506,c_out507,c_out508,c_out509,c_out510,c_out511,c_out512,c_out513,c_out514,c_out515,c_out516,c_out517,c_out518,c_out519,c_out520,c_out521,c_out522,c_out523,c_out524,c_out525,c_out526,c_out527,c_out528,c_out529,c_out530,c_out531,c_out532,c_out533,c_out534,c_out535,c_out536,c_out537,c_out538,c_out539,c_out540,c_out541,c_out542,c_out543,c_out544,c_out545,c_out546,c_out547,c_out548,c_out549,c_out550,c_out551,c_out552,c_out553,c_out554,c_out555,c_out556,c_out557,c_out558,c_out559,c_out560,c_out561,c_out562,c_out563,c_out564,c_out565,c_out566,c_out567,c_out568,c_out569,c_out570,c_out571,c_out572,c_out573,c_out574,c_out575,c_out576,c_out577,c_out578,c_out579,c_out580,c_out581,c_out582,c_out583,c_out584,c_out585,c_out586,c_out587,c_out588,c_out589,c_out590,c_out591,c_out592,c_out593,c_out594,c_out595,c_out596,c_out597,c_out598,c_out599,c_out600,c_out601,c_out602,c_out603,c_out604,c_out605,c_out606,c_out607,c_out608,c_out609,c_out610,c_out611,c_out612,c_out613,c_out614,c_out615,c_out616,c_out617,c_out618,c_out619,c_out620,c_out621,c_out622,c_out623,c_out624,c_out625,c_out626,c_out627,c_out628,c_out629,c_out630,c_out631,c_out632,c_out633,c_out634,c_out635,c_out636,c_out637,c_out638,c_out639,c_out640,c_out641,c_out642,c_out643,c_out644,c_out645,c_out646,c_out647,c_out648,c_out649,c_out650,c_out651,c_out652,c_out653,c_out654,c_out655,c_out656,c_out657,c_out658,c_out659,c_out660,c_out661,c_out662,c_out663,c_out664,c_out665,c_out666,c_out667,c_out668,c_out669,c_out670,c_out671,c_out672,c_out673,c_out674,c_out675,c_out676,c_out677,c_out678,c_out679,c_out680,c_out681,c_out682,c_out683,c_out684,c_out685,c_out686,c_out687,c_out688,c_out689,c_out690,c_out691,c_out692,c_out693,c_out694,c_out695,c_out696,c_out697,c_out698,c_out699,c_out700,c_out701,c_out702,c_out703,c_out704,c_out705,c_out706,c_out707,c_out708,c_out709,c_out710,c_out711,c_out712,c_out713,c_out714,c_out715,c_out716,c_out717,c_out718,c_out719,c_out720,c_out721,c_out722,c_out723,c_out724,c_out725,c_out726,c_out727,c_out728,c_out729,c_out730,c_out731,c_out732,c_out733,c_out734,c_out735,c_out736,c_out737,c_out738,c_out739,c_out740,c_out741,c_out742,c_out743,c_out744,c_out745,c_out746,c_out747,c_out748,c_out749,c_out750,c_out751,c_out752,c_out753,c_out754,c_out755,c_out756,c_out757,c_out758,c_out759,c_out760,c_out761,c_out762,c_out763,c_out764,c_out765,c_out766,c_out767,c_out768,c_out769,c_out770,c_out771,c_out772,c_out773,c_out774,c_out775,c_out776,c_out777,c_out778,c_out779,c_out780,c_out781,c_out782,c_out783,c_out784,c_out785,c_out786,c_out787,c_out788,c_out789,c_out790,c_out791,c_out792,c_out793,c_out794,c_out795,c_out796,c_out797,c_out798,c_out799,c_out800,c_out801,c_out802,c_out803,c_out804,c_out805,c_out806,c_out807,c_out808,c_out809,c_out810,c_out811,c_out812,c_out813,c_out814,c_out815,c_out816,c_out817,c_out818,c_out819,c_out820,c_out821,c_out822,c_out823,c_out824,c_out825,c_out826,c_out827,c_out828,c_out829,c_out830,c_out831,c_out832,c_out833,c_out834,c_out835,c_out836,c_out837,c_out838,c_out839,c_out840,c_out841,c_out842,c_out843,c_out844,c_out845,c_out846,c_out847,c_out848,c_out849,c_out850,c_out851,c_out852,c_out853,c_out854,c_out855,c_out856,c_out857,c_out858,c_out859,c_out860,c_out861,c_out862,c_out863,c_out864,c_out865,c_out866,c_out867,c_out868,c_out869,c_out870,c_out871,c_out872,c_out873,c_out874,c_out875,c_out876,c_out877,c_out878,c_out879,c_out880,c_out881,c_out882,c_out883,c_out884,c_out885,c_out886,c_out887,c_out888,c_out889,c_out890,c_out891,c_out892,c_out893,c_out894,c_out895,c_out896,c_out897,c_out898,c_out899,c_out900,c_out901,c_out902,c_out903,c_out904,c_out905,c_out906,c_out907,c_out908,c_out909,c_out910,c_out911,c_out912,c_out913,c_out914,c_out915,c_out916,c_out917,c_out918,c_out919,c_out920,c_out921,c_out922,c_out923,c_out924,c_out925,c_out926,c_out927,c_out928,c_out929,c_out930,c_out931,c_out932,c_out933,c_out934,c_out935,c_out936,c_out937,c_out938,c_out939,c_out940,c_out941,c_out942,c_out943,c_out944,c_out945,c_out946,c_out947,c_out948,c_out949,c_out950,c_out951,c_out952,c_out953,c_out954,c_out955,c_out956,c_out957,c_out958,c_out959,c_out960,c_out961,c_out962,c_out963,c_out964,c_out965,c_out966,c_out967,c_out968,c_out969,c_out970,c_out971,c_out972,c_out973,c_out974,c_out975,c_out976,c_out977,c_out978,c_out979,c_out980,c_out981,c_out982,c_out983,c_out984,c_out985,c_out986,c_out987,c_out988,c_out989,c_out990,c_out991,c_out992,c_out993,c_out994,c_out995,c_out996,c_out997,c_out998,c_out999,c_out1000,c_out1001,c_out1002,c_out1003,c_out1004,c_out1005,c_out1006,c_out1007,c_out1008,c_out1009,c_out1010,c_out1011,c_out1012,c_out1013,c_out1014,c_out1015,c_out1016,c_out1017,c_out1018,c_out1019,c_out1020,c_out1021,c_out1022,c_out1023,c_out1024,c_out1025,c_out1026,c_out1027,c_out1028,c_out1029,c_out1030,c_out1031,c_out1032,c_out1033,c_out1034,c_out1035,c_out1036,c_out1037,c_out1038,c_out1039,c_out1040,c_out1041,c_out1042,c_out1043,c_out1044,c_out1045,c_out1046,c_out1047,c_out1048,c_out1049,c_out1050,c_out1051,c_out1052,c_out1053,c_out1054,c_out1055,c_out1056,c_out1057,c_out1058,c_out1059,c_out1060,c_out1061,c_out1062,c_out1063,c_out1064,c_out1065 ,c_out1066,c_out1067,c_out1068,c_out1069,c_out1070,c_out1071,c_out1072,c_out1073,c_out1074,c_out1075,c_out1076,c_out1077,c_out1078,c_out1079,c_out1080,c_out1081,c_out1082,c_out1083 ,c_out1084,c_out1085 ,c_out1086,c_out1087,c_out1088,c_out1089,c_out1090,c_out1091,c_out1092,c_out1093,c_out1094,c_out1095,c_out1096,c_out1097,c_out1098,c_out1099,c_out1100,c_out1101,c_out1102,c_out1103,c_out1104,c_out1105,c_out1106,c_out1107,c_out1108,c_out1109,c_out1110,c_out1111,c_out1112,c_out1113,c_out1114,c_out1115,c_out1116,c_out1117,c_out1118,c_out1119,c_out1120,c_out1121,c_out1122,c_out1123,c_out1124,c_out1125,c_out1126,c_out1127,c_out1128,c_out1129,c_out1130,c_out1131,c_out1132,c_out1133,c_out1134,c_out1135,c_out1136,c_out1137,c_out1138,c_out1139,c_out1140,c_out1141,c_out1142,c_out1143,c_out1144,c_out1145,c_out1146,c_out1147,c_out1148,c_out1149,c_out1150,c_out1151,c_out1152,c_out1153,c_out1154,c_out1155,c_out1156,c_out1157,c_out1158,c_out1159,c_out1160,c_out1161,c_out1162,c_out1163,c_out1164,c_out1165,c_out1166,c_out1167,c_out1168,c_out1169,c_out1170,c_out1171,c_out1172,c_out1173,c_out1174,c_out1175,c_out1176,c_out1177,c_out1178,c_out1179,c_out1180,c_out1181,c_out1182,c_out1183,c_out1184,c_out1185,c_out1186,c_out1187,c_out1188,c_out1189,c_out1190,c_out1191,c_out1192,c_out1193,c_out1194,c_out1195,c_out1196,c_out1197,c_out1198,c_out1199,c_out1200,c_out1201,c_out1202,c_out1203,c_out1204,c_out1205,c_out1206,c_out1207,c_out1208,c_out1209,c_out1210,c_out1211,c_out1212,c_out1213,c_out1214,c_out1215,c_out1216,c_out1217,c_out1218,c_out1219,c_out1220,c_out1221,c_out1222,c_out1223,c_out1224,c_out1225,c_out1226,c_out1227,c_out1228,c_out1229,c_out1230,c_out1231,c_out1232,c_out1233,c_out1234,c_out1235,c_out1236,c_out1237,c_out1238,c_out1239,c_out1240,c_out1241,c_out1242,c_out1243,c_out1244,c_out1245,c_out1246,c_out1247,c_out1248,c_out1249,c_out1250,c_out1251,c_out1252,c_out1253,c_out1254,c_out1255,c_out1256,c_out1257,c_out1258,c_out1259,c_out1260,c_out1261,c_out1262,c_out1263,c_out1264,c_out1265,c_out1266,c_out1267,c_out1268,c_out1269,c_out1270,c_out1271,c_out1272,c_out1273,c_out1274,c_out1275,c_out1276,c_out1277,c_out1278,c_out1279,c_out1280,c_out1281,c_out1282,c_out1283,c_out1284,c_out1285,c_out1286,c_out1287,c_out1288,c_out1289,c_out1290,c_out1291,c_out1292,c_out1293,c_out1294,c_out1295,c_out1296,c_out1297,c_out1298,c_out1299,c_out1300,c_out1301,c_out1302,c_out1303,c_out1304,c_out1305,c_out1306,c_out1307,c_out1308,c_out1309,c_out1310,c_out1311,c_out1312,c_out1313,c_out1314,c_out1315,c_out1316,c_out1317,c_out1318,c_out1319,c_out1320,c_out1321,c_out1322,c_out1323,c_out1324,c_out1325,c_out1326,c_out1327,c_out1328,c_out1329,c_out1330,c_out1331,c_out1332,c_out1333,c_out1334,c_out1335,c_out1336,c_out1337,c_out1338,c_out1339,c_out1340,c_out1341,c_out1342,c_out1343,c_out1344,c_out1345,c_out1346,c_out1347,c_out1348,c_out1349,c_out1350,c_out1351,c_out1352,c_out1353,c_out1354,c_out1355,c_out1356,c_out1357,c_out1358,c_out1359,c_out1360,c_out1361,c_out1362,c_out1363,c_out1364,c_out1365,c_out1366,c_out1367,c_out1368,c_out1369,c_out1370,c_out1371,c_out1372,c_out1373,c_out1374,c_out1375,c_out1376,c_out1377,c_out1378,c_out1379,c_out1380,c_out1381,c_out1382,c_out1383,c_out1384,c_out1385,c_out1386,c_out1387,c_out1388,c_out1389,c_out1390,c_out1391,c_out1392,c_out1393,c_out1394,c_out1395,c_out1396,c_out1397,c_out1398,c_out1399,c_out1400,c_out1401,c_out1402,c_out1403,c_out1404,c_out1405,c_out1406,c_out1407,c_out1408,c_out1409,c_out1410,c_out1411,c_out1412,c_out1413,c_out1414,c_out1415,c_out1416,c_out1417,c_out1418,c_out1419,c_out1420,c_out1421,c_out1422,c_out1423,c_out1424,c_out1425,c_out1426,c_out1427,c_out1428,c_out1429,c_out1430,c_out1431,c_out1432,c_out1433,c_out1434,c_out1435,c_out1436,c_out1437,c_out1438,c_out1439,c_out1440,c_out1441,c_out1442,c_out1443,c_out1444,c_out1445,c_out1446,c_out1447,c_out1448,c_out1449,c_out1450,c_out1451,c_out1452,c_out1453,c_out1454,c_out1455,c_out1456,c_out1457,c_out1458,c_out1459,c_out1460,c_out1461,c_out1462,c_out1463,c_out1464,c_out1465,c_out1466,c_out1467,c_out1468,c_out1469,c_out1470,c_out1471,c_out1472,c_out1473,c_out1474,c_out1475,c_out1476,c_out1477,c_out1478,c_out1479,c_out1480,c_out1481,c_out1482,c_out1483,c_out1484,c_out1485,c_out1486,c_out1487,c_out1488,c_out1489,c_out1490,c_out1491,c_out1492,c_out1493,c_out1494,c_out1495,c_out1496,c_out1497,c_out1498,c_out1499,c_out1500,c_out1501,c_out1502,c_out1503,c_out1504,c_out1505,c_out1506,c_out1507,c_out1508,c_out1509,c_out1510,c_out1511,c_out1512,c_out1513,c_out1514,c_out1515,c_out1516,c_out1517,c_out1518,c_out1519,c_out1520,c_out1521,c_out1522,c_out1523,c_out1524,c_out1525,c_out1526,c_out1527,c_out1528,c_out1529,c_out1530,c_out1531,c_out1532,c_out1533,c_out1534,c_out1535,c_out1536,c_out1537,c_out1538,c_out1539,c_out1540,c_out1541,c_out1542,c_out1543,c_out1544,c_out1545,c_out1546,c_out1547,c_out1548,c_out1549,c_out1550,c_out1551,c_out1552,c_out1553,c_out1554,c_out1555,c_out1556,c_out1557,c_out1558,c_out1559,c_out1560,c_out1561,c_out1562,c_out1563,c_out1564,c_out1565,c_out1566,c_out1567,c_out1568,c_out1569,c_out1570,c_out1571,c_out1572,c_out1573,c_out1574,c_out1575,c_out1576,c_out1577,c_out1578,c_out1579,c_out1580,c_out1581,c_out1582,c_out1583,c_out1584,c_out1585,c_out1586,c_out1587,c_out1588,c_out1589,c_out1590,c_out1591,c_out1592,c_out1593,c_out1594,c_out1595,c_out1596,c_out1597,c_out1598,c_out1599,c_out1600,c_out1601,c_out1602,c_out1603,c_out1604,c_out1605,c_out1606,c_out1607,c_out1608,c_out1609,c_out1610,c_out1611,c_out1612,c_out1613,c_out1614,c_out1615,c_out1616,c_out1617,c_out1618,c_out1619,c_out1620,c_out1621,c_out1622,c_out1623,c_out1624,c_out1625,c_out1626,c_out1627,c_out1628,c_out1629,c_out1630,c_out1631,c_out1632,c_out1633,c_out1634,c_out1635,c_out1636,c_out1637,c_out1638,c_out1639,c_out1640,c_out1641,c_out1642,c_out1643,c_out1644,c_out1645,c_out1646,c_out1647,c_out1648,c_out1649,c_out1650,c_out1651,c_out1652,c_out1653,c_out1654,c_out1655,c_out1656,c_out1657,c_out1658,c_out1659,c_out1660,c_out1661,c_out1662,c_out1663,c_out1664,c_out1665,c_out1666,c_out1667,c_out1668,c_out1669,c_out1670,c_out1671,c_out1672,c_out1673,c_out1674,c_out1675,c_out1676,c_out1677,c_out1678,c_out1679,c_out1680,c_out1681,c_out1682,c_out1683,c_out1684,c_out1685,c_out1686,c_out1687,c_out1688,c_out1689,c_out1690,c_out1691,c_out1692,c_out1693,c_out1694,c_out1695,c_out1696,c_out1697,c_out1698,c_out1699,c_out1700,c_out1701,c_out1702,c_out1703,c_out1704,c_out1705,c_out1706,c_out1707,c_out1708,c_out1709,c_out1710,c_out1711,c_out1712,c_out1713,c_out1714,c_out1715,c_out1716,c_out1717,c_out1718,c_out1719,c_out1720,c_out1721,c_out1722,c_out1723,c_out1724,c_out1725,c_out1726,c_out1727,c_out1728,c_out1729,c_out1730,c_out1731,c_out1732,c_out1733,c_out1734,c_out1735,c_out1736,c_out1737,c_out1738,c_out1739,c_out1740,c_out1741,c_out1742,c_out1743,c_out1744,c_out1745,c_out1746,c_out1747,c_out1748,c_out1749,c_out1750,c_out1751,c_out1752,c_out1753,c_out1754,c_out1755,c_out1756,c_out1757,c_out1758,c_out1759,c_out1760,c_out1761,c_out1762,c_out1763,c_out1764,c_out1765,c_out1766,c_out1767,c_out1768,c_out1769,c_out1770,c_out1771,c_out1772,c_out1773,c_out1774,c_out1775,c_out1776,c_out1777,c_out1778,c_out1779,c_out1780,c_out1781,c_out1782,c_out1783,c_out1784,c_out1785,c_out1786,c_out1787,c_out1788,c_out1789,c_out1790,c_out1791,c_out1792,c_out1793,c_out1794,c_out1795,c_out1796,c_out1797,c_out1798,c_out1799,c_out1800,c_out1801,c_out1802,c_out1803,c_out1804,c_out1805,c_out1806,c_out1807,c_out1808,c_out1809,c_out1810,c_out1811,c_out1812,c_out1813,c_out1814,c_out1815,c_out1816,c_out1817,c_out1818,c_out1819,c_out1820,c_out1821,c_out1822,c_out1823,c_out1824,c_out1825,c_out1826,c_out1827,c_out1828,c_out1829,c_out1830,c_out1831,c_out1832,c_out1833,c_out1834,c_out1835,c_out1836,c_out1837,c_out1838,c_out1839,c_out1840,c_out1841,c_out1842,c_out1843,c_out1844,c_out1845,c_out1846,c_out1847,c_out1848,c_out1849,c_out1850,c_out1851,c_out1852,c_out1853,c_out1854,c_out1855,c_out1856,c_out1857,c_out1858,c_out1859,c_out1860,c_out1861,c_out1862,c_out1863,c_out1864,c_out1865,c_out1866,c_out1867,c_out1868,c_out1869,c_out1870,c_out1871,c_out1872,c_out1873,c_out1874,c_out1875,c_out1876,c_out1877,c_out1878,c_out1879,c_out1880,c_out1881,c_out1882,c_out1883,c_out1884,c_out1885,c_out1886,c_out1887,c_out1888,c_out1889,c_out1890,c_out1891,c_out1892,c_out1893,c_out1894,c_out1895,c_out1896,c_out1897,c_out1898,c_out1899,c_out1900,c_out1901,c_out1902,c_out1903,c_out1904,c_out1905,c_out1906,c_out1907,c_out1908,c_out1909,c_out1910,c_out1911,c_out1912,c_out1913,c_out1914,c_out1915,c_out1916,c_out1917,c_out1918,c_out1919,c_out1920,c_out1921,c_out1922,c_out1923,c_out1924,c_out1925,c_out1926,c_out1927,c_out1928,c_out1929,c_out1930,c_out1931,c_out1932,c_out1933,c_out1934,c_out1935,c_out1936,c_out1937,c_out1938,c_out1939,c_out1940,c_out1941,c_out1942,c_out1943,c_out1944,c_out1945,c_out1946,c_out1947,c_out1948,c_out1949,c_out1950,c_out1951,c_out1952,c_out1953,c_out1954,c_out1955,c_out1956,c_out1957,c_out1958,c_out1959,c_out1960,c_out1961,c_out1962,c_out1963,c_out1964,c_out1965,c_out1966,c_out1967,c_out1968,c_out1969,c_out1970,c_out1971,c_out1972,c_out1973,c_out1974,c_out1975,c_out1976,c_out1977,c_out1978,c_out1979,c_out1980,c_out1981,c_out1982,c_out1983,c_out1984,c_out1985,c_out1986,c_out1987,c_out1988,c_out1989,c_out1990,c_out1991,c_out1992,c_out1993,c_out1994,c_out1995,c_out1996,c_out1997,c_out1998,c_out1999,c_out2000,c_out2001,c_out2002,c_out2003,c_out2004,c_out2005,c_out2006,c_out2007,c_out2008,c_out2009,c_out2010,c_out2011,c_out2012,c_out2013,c_out2014,c_out2015,c_out2016,c_out2017,c_out2018,c_out2019,c_out2020,c_out2021,c_out2022,c_out2023,c_out2024,c_out2025,c_out2026,c_out2027,c_out2028,c_out2029,c_out2030,c_out2031,c_out2032,c_out2033,c_out2034,c_out2035,c_out2036,c_out2037,c_out2038,c_out2039,c_out2040,c_out2041,c_out2042,c_out2043,c_out2044,c_out2045,c_out2046,c_out2047,out_act,out_weight);

parameter WIDTH = 8;
parameter C_WIDTH = 32;

input clk,rstn;
input [256*WIDTH-1:0] activation;
input [256*WIDTH-1:0] weight;
input control;
output [32*C_WIDTH-1:0] c_out0;
output [32*C_WIDTH-1:0] c_out1;
output [32*C_WIDTH-1:0] c_out2;
output [32*C_WIDTH-1:0] c_out3;
output [32*C_WIDTH-1:0] c_out4;
output [32*C_WIDTH-1:0] c_out5;
output [32*C_WIDTH-1:0] c_out6;
output [32*C_WIDTH-1:0] c_out7;
output [32*C_WIDTH-1:0] c_out8;
output [32*C_WIDTH-1:0] c_out9;
output [32*C_WIDTH-1:0] c_out10;
output [32*C_WIDTH-1:0] c_out11;
output [32*C_WIDTH-1:0] c_out12;
output [32*C_WIDTH-1:0] c_out13;
output [32*C_WIDTH-1:0] c_out14;
output [32*C_WIDTH-1:0] c_out15;
output [32*C_WIDTH-1:0] c_out16;
output [32*C_WIDTH-1:0] c_out17;
output [32*C_WIDTH-1:0] c_out18;
output [32*C_WIDTH-1:0] c_out19;
output [32*C_WIDTH-1:0] c_out20;
output [32*C_WIDTH-1:0] c_out21;
output [32*C_WIDTH-1:0] c_out22;
output [32*C_WIDTH-1:0] c_out23;
output [32*C_WIDTH-1:0] c_out24;
output [32*C_WIDTH-1:0] c_out25;
output [32*C_WIDTH-1:0] c_out26;
output [32*C_WIDTH-1:0] c_out27;
output [32*C_WIDTH-1:0] c_out28;
output [32*C_WIDTH-1:0] c_out29;
output [32*C_WIDTH-1:0] c_out30;
output [32*C_WIDTH-1:0] c_out31;
output [32*C_WIDTH-1:0] c_out32;
output [32*C_WIDTH-1:0] c_out33;
output [32*C_WIDTH-1:0] c_out34;
output [32*C_WIDTH-1:0] c_out35;
output [32*C_WIDTH-1:0] c_out36;
output [32*C_WIDTH-1:0] c_out37;
output [32*C_WIDTH-1:0] c_out38;
output [32*C_WIDTH-1:0] c_out39;
output [32*C_WIDTH-1:0] c_out40;
output [32*C_WIDTH-1:0] c_out41;
output [32*C_WIDTH-1:0] c_out42;
output [32*C_WIDTH-1:0] c_out43;
output [32*C_WIDTH-1:0] c_out44;
output [32*C_WIDTH-1:0] c_out45;
output [32*C_WIDTH-1:0] c_out46;
output [32*C_WIDTH-1:0] c_out47;
output [32*C_WIDTH-1:0] c_out48;
output [32*C_WIDTH-1:0] c_out49;
output [32*C_WIDTH-1:0] c_out50;
output [32*C_WIDTH-1:0] c_out51;
output [32*C_WIDTH-1:0] c_out52;
output [32*C_WIDTH-1:0] c_out53;
output [32*C_WIDTH-1:0] c_out54;
output [32*C_WIDTH-1:0] c_out55;
output [32*C_WIDTH-1:0] c_out56;
output [32*C_WIDTH-1:0] c_out57;
output [32*C_WIDTH-1:0] c_out58;
output [32*C_WIDTH-1:0] c_out59;
output [32*C_WIDTH-1:0] c_out60;
output [32*C_WIDTH-1:0] c_out61;
output [32*C_WIDTH-1:0] c_out62;
output [32*C_WIDTH-1:0] c_out63;
output [32*C_WIDTH-1:0] c_out64;
output [32*C_WIDTH-1:0] c_out65;
output [32*C_WIDTH-1:0] c_out66;
output [32*C_WIDTH-1:0] c_out67;
output [32*C_WIDTH-1:0] c_out68;
output [32*C_WIDTH-1:0] c_out69;
output [32*C_WIDTH-1:0] c_out70;
output [32*C_WIDTH-1:0] c_out71;
output [32*C_WIDTH-1:0] c_out72;
output [32*C_WIDTH-1:0] c_out73;
output [32*C_WIDTH-1:0] c_out74;
output [32*C_WIDTH-1:0] c_out75;
output [32*C_WIDTH-1:0] c_out76;
output [32*C_WIDTH-1:0] c_out77;
output [32*C_WIDTH-1:0] c_out78;
output [32*C_WIDTH-1:0] c_out79;
output [32*C_WIDTH-1:0] c_out80;
output [32*C_WIDTH-1:0] c_out81;
output [32*C_WIDTH-1:0] c_out82;
output [32*C_WIDTH-1:0] c_out83;
output [32*C_WIDTH-1:0] c_out84;
output [32*C_WIDTH-1:0] c_out85;
output [32*C_WIDTH-1:0] c_out86;
output [32*C_WIDTH-1:0] c_out87;
output [32*C_WIDTH-1:0] c_out88;
output [32*C_WIDTH-1:0] c_out89;
output [32*C_WIDTH-1:0] c_out90;
output [32*C_WIDTH-1:0] c_out91;
output [32*C_WIDTH-1:0] c_out92;
output [32*C_WIDTH-1:0] c_out93;
output [32*C_WIDTH-1:0] c_out94;
output [32*C_WIDTH-1:0] c_out95;
output [32*C_WIDTH-1:0] c_out96;
output [32*C_WIDTH-1:0] c_out97;
output [32*C_WIDTH-1:0] c_out98;
output [32*C_WIDTH-1:0] c_out99;
output [32*C_WIDTH-1:0] c_out100;
output [32*C_WIDTH-1:0] c_out101;
output [32*C_WIDTH-1:0] c_out102;
output [32*C_WIDTH-1:0] c_out103;
output [32*C_WIDTH-1:0] c_out104;
output [32*C_WIDTH-1:0] c_out105;
output [32*C_WIDTH-1:0] c_out106;
output [32*C_WIDTH-1:0] c_out107;
output [32*C_WIDTH-1:0] c_out108;
output [32*C_WIDTH-1:0] c_out109;
output [32*C_WIDTH-1:0] c_out110;
output [32*C_WIDTH-1:0] c_out111;
output [32*C_WIDTH-1:0] c_out112;
output [32*C_WIDTH-1:0] c_out113;
output [32*C_WIDTH-1:0] c_out114;
output [32*C_WIDTH-1:0] c_out115;
output [32*C_WIDTH-1:0] c_out116;
output [32*C_WIDTH-1:0] c_out117;
output [32*C_WIDTH-1:0] c_out118;
output [32*C_WIDTH-1:0] c_out119;
output [32*C_WIDTH-1:0] c_out120;
output [32*C_WIDTH-1:0] c_out121;
output [32*C_WIDTH-1:0] c_out122;
output [32*C_WIDTH-1:0] c_out123;
output [32*C_WIDTH-1:0] c_out124;
output [32*C_WIDTH-1:0] c_out125;
output [32*C_WIDTH-1:0] c_out126;
output [32*C_WIDTH-1:0] c_out127;
output [32*C_WIDTH-1:0] c_out128;
output [32*C_WIDTH-1:0] c_out129;
output [32*C_WIDTH-1:0] c_out130;
output [32*C_WIDTH-1:0] c_out131;
output [32*C_WIDTH-1:0] c_out132;
output [32*C_WIDTH-1:0] c_out133;
output [32*C_WIDTH-1:0] c_out134;
output [32*C_WIDTH-1:0] c_out135;
output [32*C_WIDTH-1:0] c_out136;
output [32*C_WIDTH-1:0] c_out137;
output [32*C_WIDTH-1:0] c_out138;
output [32*C_WIDTH-1:0] c_out139;
output [32*C_WIDTH-1:0] c_out140;
output [32*C_WIDTH-1:0] c_out141;
output [32*C_WIDTH-1:0] c_out142;
output [32*C_WIDTH-1:0] c_out143;
output [32*C_WIDTH-1:0] c_out144;
output [32*C_WIDTH-1:0] c_out145;
output [32*C_WIDTH-1:0] c_out146;
output [32*C_WIDTH-1:0] c_out147;
output [32*C_WIDTH-1:0] c_out148;
output [32*C_WIDTH-1:0] c_out149;
output [32*C_WIDTH-1:0] c_out150;
output [32*C_WIDTH-1:0] c_out151;
output [32*C_WIDTH-1:0] c_out152;
output [32*C_WIDTH-1:0] c_out153;
output [32*C_WIDTH-1:0] c_out154;
output [32*C_WIDTH-1:0] c_out155;
output [32*C_WIDTH-1:0] c_out156;
output [32*C_WIDTH-1:0] c_out157;
output [32*C_WIDTH-1:0] c_out158;
output [32*C_WIDTH-1:0] c_out159;
output [32*C_WIDTH-1:0] c_out160;
output [32*C_WIDTH-1:0] c_out161;
output [32*C_WIDTH-1:0] c_out162;
output [32*C_WIDTH-1:0] c_out163;
output [32*C_WIDTH-1:0] c_out164;
output [32*C_WIDTH-1:0] c_out165;
output [32*C_WIDTH-1:0] c_out166;
output [32*C_WIDTH-1:0] c_out167;
output [32*C_WIDTH-1:0] c_out168;
output [32*C_WIDTH-1:0] c_out169;
output [32*C_WIDTH-1:0] c_out170;
output [32*C_WIDTH-1:0] c_out171;
output [32*C_WIDTH-1:0] c_out172;
output [32*C_WIDTH-1:0] c_out173;
output [32*C_WIDTH-1:0] c_out174;
output [32*C_WIDTH-1:0] c_out175;
output [32*C_WIDTH-1:0] c_out176;
output [32*C_WIDTH-1:0] c_out177;
output [32*C_WIDTH-1:0] c_out178;
output [32*C_WIDTH-1:0] c_out179;
output [32*C_WIDTH-1:0] c_out180;
output [32*C_WIDTH-1:0] c_out181;
output [32*C_WIDTH-1:0] c_out182;
output [32*C_WIDTH-1:0] c_out183;
output [32*C_WIDTH-1:0] c_out184;
output [32*C_WIDTH-1:0] c_out185;
output [32*C_WIDTH-1:0] c_out186;
output [32*C_WIDTH-1:0] c_out187;
output [32*C_WIDTH-1:0] c_out188;
output [32*C_WIDTH-1:0] c_out189;
output [32*C_WIDTH-1:0] c_out190;
output [32*C_WIDTH-1:0] c_out191;
output [32*C_WIDTH-1:0] c_out192;
output [32*C_WIDTH-1:0] c_out193;
output [32*C_WIDTH-1:0] c_out194;
output [32*C_WIDTH-1:0] c_out195;
output [32*C_WIDTH-1:0] c_out196;
output [32*C_WIDTH-1:0] c_out197;
output [32*C_WIDTH-1:0] c_out198;
output [32*C_WIDTH-1:0] c_out199;
output [32*C_WIDTH-1:0] c_out200;
output [32*C_WIDTH-1:0] c_out201;
output [32*C_WIDTH-1:0] c_out202;
output [32*C_WIDTH-1:0] c_out203;
output [32*C_WIDTH-1:0] c_out204;
output [32*C_WIDTH-1:0] c_out205;
output [32*C_WIDTH-1:0] c_out206;
output [32*C_WIDTH-1:0] c_out207;
output [32*C_WIDTH-1:0] c_out208;
output [32*C_WIDTH-1:0] c_out209;
output [32*C_WIDTH-1:0] c_out210;
output [32*C_WIDTH-1:0] c_out211;
output [32*C_WIDTH-1:0] c_out212;
output [32*C_WIDTH-1:0] c_out213;
output [32*C_WIDTH-1:0] c_out214;
output [32*C_WIDTH-1:0] c_out215;
output [32*C_WIDTH-1:0] c_out216;
output [32*C_WIDTH-1:0] c_out217;
output [32*C_WIDTH-1:0] c_out218;
output [32*C_WIDTH-1:0] c_out219;
output [32*C_WIDTH-1:0] c_out220;
output [32*C_WIDTH-1:0] c_out221;
output [32*C_WIDTH-1:0] c_out222;
output [32*C_WIDTH-1:0] c_out223;
output [32*C_WIDTH-1:0] c_out224;
output [32*C_WIDTH-1:0] c_out225;
output [32*C_WIDTH-1:0] c_out226;
output [32*C_WIDTH-1:0] c_out227;
output [32*C_WIDTH-1:0] c_out228;
output [32*C_WIDTH-1:0] c_out229;
output [32*C_WIDTH-1:0] c_out230;
output [32*C_WIDTH-1:0] c_out231;
output [32*C_WIDTH-1:0] c_out232;
output [32*C_WIDTH-1:0] c_out233;
output [32*C_WIDTH-1:0] c_out234;
output [32*C_WIDTH-1:0] c_out235;
output [32*C_WIDTH-1:0] c_out236;
output [32*C_WIDTH-1:0] c_out237;
output [32*C_WIDTH-1:0] c_out238;
output [32*C_WIDTH-1:0] c_out239;
output [32*C_WIDTH-1:0] c_out240;
output [32*C_WIDTH-1:0] c_out241;
output [32*C_WIDTH-1:0] c_out242;
output [32*C_WIDTH-1:0] c_out243;
output [32*C_WIDTH-1:0] c_out244;
output [32*C_WIDTH-1:0] c_out245;
output [32*C_WIDTH-1:0] c_out246;
output [32*C_WIDTH-1:0] c_out247;
output [32*C_WIDTH-1:0] c_out248;
output [32*C_WIDTH-1:0] c_out249;
output [32*C_WIDTH-1:0] c_out250;
output [32*C_WIDTH-1:0] c_out251;
output [32*C_WIDTH-1:0] c_out252;
output [32*C_WIDTH-1:0] c_out253;
output [32*C_WIDTH-1:0] c_out254;
output [32*C_WIDTH-1:0] c_out255;
output [32*C_WIDTH-1:0] c_out256;
output [32*C_WIDTH-1:0] c_out257;
output [32*C_WIDTH-1:0] c_out258;
output [32*C_WIDTH-1:0] c_out259;
output [32*C_WIDTH-1:0] c_out260;
output [32*C_WIDTH-1:0] c_out261;
output [32*C_WIDTH-1:0] c_out262;
output [32*C_WIDTH-1:0] c_out263;
output [32*C_WIDTH-1:0] c_out264;
output [32*C_WIDTH-1:0] c_out265;
output [32*C_WIDTH-1:0] c_out266;
output [32*C_WIDTH-1:0] c_out267;
output [32*C_WIDTH-1:0] c_out268;
output [32*C_WIDTH-1:0] c_out269;
output [32*C_WIDTH-1:0] c_out270;
output [32*C_WIDTH-1:0] c_out271;
output [32*C_WIDTH-1:0] c_out272;
output [32*C_WIDTH-1:0] c_out273;
output [32*C_WIDTH-1:0] c_out274;
output [32*C_WIDTH-1:0] c_out275;
output [32*C_WIDTH-1:0] c_out276;
output [32*C_WIDTH-1:0] c_out277;
output [32*C_WIDTH-1:0] c_out278;
output [32*C_WIDTH-1:0] c_out279;
output [32*C_WIDTH-1:0] c_out280;
output [32*C_WIDTH-1:0] c_out281;
output [32*C_WIDTH-1:0] c_out282;
output [32*C_WIDTH-1:0] c_out283;
output [32*C_WIDTH-1:0] c_out284;
output [32*C_WIDTH-1:0] c_out285;
output [32*C_WIDTH-1:0] c_out286;
output [32*C_WIDTH-1:0] c_out287;
output [32*C_WIDTH-1:0] c_out288;
output [32*C_WIDTH-1:0] c_out289;
output [32*C_WIDTH-1:0] c_out290;
output [32*C_WIDTH-1:0] c_out291;
output [32*C_WIDTH-1:0] c_out292;
output [32*C_WIDTH-1:0] c_out293;
output [32*C_WIDTH-1:0] c_out294;
output [32*C_WIDTH-1:0] c_out295;
output [32*C_WIDTH-1:0] c_out296;
output [32*C_WIDTH-1:0] c_out297;
output [32*C_WIDTH-1:0] c_out298;
output [32*C_WIDTH-1:0] c_out299;
output [32*C_WIDTH-1:0] c_out300;
output [32*C_WIDTH-1:0] c_out301;
output [32*C_WIDTH-1:0] c_out302;
output [32*C_WIDTH-1:0] c_out303;
output [32*C_WIDTH-1:0] c_out304;
output [32*C_WIDTH-1:0] c_out305;
output [32*C_WIDTH-1:0] c_out306;
output [32*C_WIDTH-1:0] c_out307;
output [32*C_WIDTH-1:0] c_out308;
output [32*C_WIDTH-1:0] c_out309;
output [32*C_WIDTH-1:0] c_out310;
output [32*C_WIDTH-1:0] c_out311;
output [32*C_WIDTH-1:0] c_out312;
output [32*C_WIDTH-1:0] c_out313;
output [32*C_WIDTH-1:0] c_out314;
output [32*C_WIDTH-1:0] c_out315;
output [32*C_WIDTH-1:0] c_out316;
output [32*C_WIDTH-1:0] c_out317;
output [32*C_WIDTH-1:0] c_out318;
output [32*C_WIDTH-1:0] c_out319;
output [32*C_WIDTH-1:0] c_out320;
output [32*C_WIDTH-1:0] c_out321;
output [32*C_WIDTH-1:0] c_out322;
output [32*C_WIDTH-1:0] c_out323;
output [32*C_WIDTH-1:0] c_out324;
output [32*C_WIDTH-1:0] c_out325;
output [32*C_WIDTH-1:0] c_out326;
output [32*C_WIDTH-1:0] c_out327;
output [32*C_WIDTH-1:0] c_out328;
output [32*C_WIDTH-1:0] c_out329;
output [32*C_WIDTH-1:0] c_out330;
output [32*C_WIDTH-1:0] c_out331;
output [32*C_WIDTH-1:0] c_out332;
output [32*C_WIDTH-1:0] c_out333;
output [32*C_WIDTH-1:0] c_out334;
output [32*C_WIDTH-1:0] c_out335;
output [32*C_WIDTH-1:0] c_out336;
output [32*C_WIDTH-1:0] c_out337;
output [32*C_WIDTH-1:0] c_out338;
output [32*C_WIDTH-1:0] c_out339;
output [32*C_WIDTH-1:0] c_out340;
output [32*C_WIDTH-1:0] c_out341;
output [32*C_WIDTH-1:0] c_out342;
output [32*C_WIDTH-1:0] c_out343;
output [32*C_WIDTH-1:0] c_out344;
output [32*C_WIDTH-1:0] c_out345;
output [32*C_WIDTH-1:0] c_out346;
output [32*C_WIDTH-1:0] c_out347;
output [32*C_WIDTH-1:0] c_out348;
output [32*C_WIDTH-1:0] c_out349;
output [32*C_WIDTH-1:0] c_out350;
output [32*C_WIDTH-1:0] c_out351;
output [32*C_WIDTH-1:0] c_out352;
output [32*C_WIDTH-1:0] c_out353;
output [32*C_WIDTH-1:0] c_out354;
output [32*C_WIDTH-1:0] c_out355;
output [32*C_WIDTH-1:0] c_out356;
output [32*C_WIDTH-1:0] c_out357;
output [32*C_WIDTH-1:0] c_out358;
output [32*C_WIDTH-1:0] c_out359;
output [32*C_WIDTH-1:0] c_out360;
output [32*C_WIDTH-1:0] c_out361;
output [32*C_WIDTH-1:0] c_out362;
output [32*C_WIDTH-1:0] c_out363;
output [32*C_WIDTH-1:0] c_out364;
output [32*C_WIDTH-1:0] c_out365;
output [32*C_WIDTH-1:0] c_out366;
output [32*C_WIDTH-1:0] c_out367;
output [32*C_WIDTH-1:0] c_out368;
output [32*C_WIDTH-1:0] c_out369;
output [32*C_WIDTH-1:0] c_out370;
output [32*C_WIDTH-1:0] c_out371;
output [32*C_WIDTH-1:0] c_out372;
output [32*C_WIDTH-1:0] c_out373;
output [32*C_WIDTH-1:0] c_out374;
output [32*C_WIDTH-1:0] c_out375;
output [32*C_WIDTH-1:0] c_out376;
output [32*C_WIDTH-1:0] c_out377;
output [32*C_WIDTH-1:0] c_out378;
output [32*C_WIDTH-1:0] c_out379;
output [32*C_WIDTH-1:0] c_out380;
output [32*C_WIDTH-1:0] c_out381;
output [32*C_WIDTH-1:0] c_out382;
output [32*C_WIDTH-1:0] c_out383;
output [32*C_WIDTH-1:0] c_out384;
output [32*C_WIDTH-1:0] c_out385;
output [32*C_WIDTH-1:0] c_out386;
output [32*C_WIDTH-1:0] c_out387;
output [32*C_WIDTH-1:0] c_out388;
output [32*C_WIDTH-1:0] c_out389;
output [32*C_WIDTH-1:0] c_out390;
output [32*C_WIDTH-1:0] c_out391;
output [32*C_WIDTH-1:0] c_out392;
output [32*C_WIDTH-1:0] c_out393;
output [32*C_WIDTH-1:0] c_out394;
output [32*C_WIDTH-1:0] c_out395;
output [32*C_WIDTH-1:0] c_out396;
output [32*C_WIDTH-1:0] c_out397;
output [32*C_WIDTH-1:0] c_out398;
output [32*C_WIDTH-1:0] c_out399;
output [32*C_WIDTH-1:0] c_out400;
output [32*C_WIDTH-1:0] c_out401;
output [32*C_WIDTH-1:0] c_out402;
output [32*C_WIDTH-1:0] c_out403;
output [32*C_WIDTH-1:0] c_out404;
output [32*C_WIDTH-1:0] c_out405;
output [32*C_WIDTH-1:0] c_out406;
output [32*C_WIDTH-1:0] c_out407;
output [32*C_WIDTH-1:0] c_out408;
output [32*C_WIDTH-1:0] c_out409;
output [32*C_WIDTH-1:0] c_out410;
output [32*C_WIDTH-1:0] c_out411;
output [32*C_WIDTH-1:0] c_out412;
output [32*C_WIDTH-1:0] c_out413;
output [32*C_WIDTH-1:0] c_out414;
output [32*C_WIDTH-1:0] c_out415;
output [32*C_WIDTH-1:0] c_out416;
output [32*C_WIDTH-1:0] c_out417;
output [32*C_WIDTH-1:0] c_out418;
output [32*C_WIDTH-1:0] c_out419;
output [32*C_WIDTH-1:0] c_out420;
output [32*C_WIDTH-1:0] c_out421;
output [32*C_WIDTH-1:0] c_out422;
output [32*C_WIDTH-1:0] c_out423;
output [32*C_WIDTH-1:0] c_out424;
output [32*C_WIDTH-1:0] c_out425;
output [32*C_WIDTH-1:0] c_out426;
output [32*C_WIDTH-1:0] c_out427;
output [32*C_WIDTH-1:0] c_out428;
output [32*C_WIDTH-1:0] c_out429;
output [32*C_WIDTH-1:0] c_out430;
output [32*C_WIDTH-1:0] c_out431;
output [32*C_WIDTH-1:0] c_out432;
output [32*C_WIDTH-1:0] c_out433;
output [32*C_WIDTH-1:0] c_out434;
output [32*C_WIDTH-1:0] c_out435;
output [32*C_WIDTH-1:0] c_out436;
output [32*C_WIDTH-1:0] c_out437;
output [32*C_WIDTH-1:0] c_out438;
output [32*C_WIDTH-1:0] c_out439;
output [32*C_WIDTH-1:0] c_out440;
output [32*C_WIDTH-1:0] c_out441;
output [32*C_WIDTH-1:0] c_out442;
output [32*C_WIDTH-1:0] c_out443;
output [32*C_WIDTH-1:0] c_out444;
output [32*C_WIDTH-1:0] c_out445;
output [32*C_WIDTH-1:0] c_out446;
output [32*C_WIDTH-1:0] c_out447;
output [32*C_WIDTH-1:0] c_out448;
output [32*C_WIDTH-1:0] c_out449;
output [32*C_WIDTH-1:0] c_out450;
output [32*C_WIDTH-1:0] c_out451;
output [32*C_WIDTH-1:0] c_out452;
output [32*C_WIDTH-1:0] c_out453;
output [32*C_WIDTH-1:0] c_out454;
output [32*C_WIDTH-1:0] c_out455;
output [32*C_WIDTH-1:0] c_out456;
output [32*C_WIDTH-1:0] c_out457;
output [32*C_WIDTH-1:0] c_out458;
output [32*C_WIDTH-1:0] c_out459;
output [32*C_WIDTH-1:0] c_out460;
output [32*C_WIDTH-1:0] c_out461;
output [32*C_WIDTH-1:0] c_out462;
output [32*C_WIDTH-1:0] c_out463;
output [32*C_WIDTH-1:0] c_out464;
output [32*C_WIDTH-1:0] c_out465;
output [32*C_WIDTH-1:0] c_out466;
output [32*C_WIDTH-1:0] c_out467;
output [32*C_WIDTH-1:0] c_out468;
output [32*C_WIDTH-1:0] c_out469;
output [32*C_WIDTH-1:0] c_out470;
output [32*C_WIDTH-1:0] c_out471;
output [32*C_WIDTH-1:0] c_out472;
output [32*C_WIDTH-1:0] c_out473;
output [32*C_WIDTH-1:0] c_out474;
output [32*C_WIDTH-1:0] c_out475;
output [32*C_WIDTH-1:0] c_out476;
output [32*C_WIDTH-1:0] c_out477;
output [32*C_WIDTH-1:0] c_out478;
output [32*C_WIDTH-1:0] c_out479;
output [32*C_WIDTH-1:0] c_out480;
output [32*C_WIDTH-1:0] c_out481;
output [32*C_WIDTH-1:0] c_out482;
output [32*C_WIDTH-1:0] c_out483;
output [32*C_WIDTH-1:0] c_out484;
output [32*C_WIDTH-1:0] c_out485;
output [32*C_WIDTH-1:0] c_out486;
output [32*C_WIDTH-1:0] c_out487;
output [32*C_WIDTH-1:0] c_out488;
output [32*C_WIDTH-1:0] c_out489;
output [32*C_WIDTH-1:0] c_out490;
output [32*C_WIDTH-1:0] c_out491;
output [32*C_WIDTH-1:0] c_out492;
output [32*C_WIDTH-1:0] c_out493;
output [32*C_WIDTH-1:0] c_out494;
output [32*C_WIDTH-1:0] c_out495;
output [32*C_WIDTH-1:0] c_out496;
output [32*C_WIDTH-1:0] c_out497;
output [32*C_WIDTH-1:0] c_out498;
output [32*C_WIDTH-1:0] c_out499;
output [32*C_WIDTH-1:0] c_out500;
output [32*C_WIDTH-1:0] c_out501;
output [32*C_WIDTH-1:0] c_out502;
output [32*C_WIDTH-1:0] c_out503;
output [32*C_WIDTH-1:0] c_out504;
output [32*C_WIDTH-1:0] c_out505;
output [32*C_WIDTH-1:0] c_out506;
output [32*C_WIDTH-1:0] c_out507;
output [32*C_WIDTH-1:0] c_out508;
output [32*C_WIDTH-1:0] c_out509;
output [32*C_WIDTH-1:0] c_out510;
output [32*C_WIDTH-1:0] c_out511;
output [32*C_WIDTH-1:0] c_out512;
output [32*C_WIDTH-1:0] c_out513;
output [32*C_WIDTH-1:0] c_out514;
output [32*C_WIDTH-1:0] c_out515;
output [32*C_WIDTH-1:0] c_out516;
output [32*C_WIDTH-1:0] c_out517;
output [32*C_WIDTH-1:0] c_out518;
output [32*C_WIDTH-1:0] c_out519;
output [32*C_WIDTH-1:0] c_out520;
output [32*C_WIDTH-1:0] c_out521;
output [32*C_WIDTH-1:0] c_out522;
output [32*C_WIDTH-1:0] c_out523;
output [32*C_WIDTH-1:0] c_out524;
output [32*C_WIDTH-1:0] c_out525;
output [32*C_WIDTH-1:0] c_out526;
output [32*C_WIDTH-1:0] c_out527;
output [32*C_WIDTH-1:0] c_out528;
output [32*C_WIDTH-1:0] c_out529;
output [32*C_WIDTH-1:0] c_out530;
output [32*C_WIDTH-1:0] c_out531;
output [32*C_WIDTH-1:0] c_out532;
output [32*C_WIDTH-1:0] c_out533;
output [32*C_WIDTH-1:0] c_out534;
output [32*C_WIDTH-1:0] c_out535;
output [32*C_WIDTH-1:0] c_out536;
output [32*C_WIDTH-1:0] c_out537;
output [32*C_WIDTH-1:0] c_out538;
output [32*C_WIDTH-1:0] c_out539;
output [32*C_WIDTH-1:0] c_out540;
output [32*C_WIDTH-1:0] c_out541;
output [32*C_WIDTH-1:0] c_out542;
output [32*C_WIDTH-1:0] c_out543;
output [32*C_WIDTH-1:0] c_out544;
output [32*C_WIDTH-1:0] c_out545;
output [32*C_WIDTH-1:0] c_out546;
output [32*C_WIDTH-1:0] c_out547;
output [32*C_WIDTH-1:0] c_out548;
output [32*C_WIDTH-1:0] c_out549;
output [32*C_WIDTH-1:0] c_out550;
output [32*C_WIDTH-1:0] c_out551;
output [32*C_WIDTH-1:0] c_out552;
output [32*C_WIDTH-1:0] c_out553;
output [32*C_WIDTH-1:0] c_out554;
output [32*C_WIDTH-1:0] c_out555;
output [32*C_WIDTH-1:0] c_out556;
output [32*C_WIDTH-1:0] c_out557;
output [32*C_WIDTH-1:0] c_out558;
output [32*C_WIDTH-1:0] c_out559;
output [32*C_WIDTH-1:0] c_out560;
output [32*C_WIDTH-1:0] c_out561;
output [32*C_WIDTH-1:0] c_out562;
output [32*C_WIDTH-1:0] c_out563;
output [32*C_WIDTH-1:0] c_out564;
output [32*C_WIDTH-1:0] c_out565;
output [32*C_WIDTH-1:0] c_out566;
output [32*C_WIDTH-1:0] c_out567;
output [32*C_WIDTH-1:0] c_out568;
output [32*C_WIDTH-1:0] c_out569;
output [32*C_WIDTH-1:0] c_out570;
output [32*C_WIDTH-1:0] c_out571;
output [32*C_WIDTH-1:0] c_out572;
output [32*C_WIDTH-1:0] c_out573;
output [32*C_WIDTH-1:0] c_out574;
output [32*C_WIDTH-1:0] c_out575;
output [32*C_WIDTH-1:0] c_out576;
output [32*C_WIDTH-1:0] c_out577;
output [32*C_WIDTH-1:0] c_out578;
output [32*C_WIDTH-1:0] c_out579;
output [32*C_WIDTH-1:0] c_out580;
output [32*C_WIDTH-1:0] c_out581;
output [32*C_WIDTH-1:0] c_out582;
output [32*C_WIDTH-1:0] c_out583;
output [32*C_WIDTH-1:0] c_out584;
output [32*C_WIDTH-1:0] c_out585;
output [32*C_WIDTH-1:0] c_out586;
output [32*C_WIDTH-1:0] c_out587;
output [32*C_WIDTH-1:0] c_out588;
output [32*C_WIDTH-1:0] c_out589;
output [32*C_WIDTH-1:0] c_out590;
output [32*C_WIDTH-1:0] c_out591;
output [32*C_WIDTH-1:0] c_out592;
output [32*C_WIDTH-1:0] c_out593;
output [32*C_WIDTH-1:0] c_out594;
output [32*C_WIDTH-1:0] c_out595;
output [32*C_WIDTH-1:0] c_out596;
output [32*C_WIDTH-1:0] c_out597;
output [32*C_WIDTH-1:0] c_out598;
output [32*C_WIDTH-1:0] c_out599;
output [32*C_WIDTH-1:0] c_out600;
output [32*C_WIDTH-1:0] c_out601;
output [32*C_WIDTH-1:0] c_out602;
output [32*C_WIDTH-1:0] c_out603;
output [32*C_WIDTH-1:0] c_out604;
output [32*C_WIDTH-1:0] c_out605;
output [32*C_WIDTH-1:0] c_out606;
output [32*C_WIDTH-1:0] c_out607;
output [32*C_WIDTH-1:0] c_out608;
output [32*C_WIDTH-1:0] c_out609;
output [32*C_WIDTH-1:0] c_out610;
output [32*C_WIDTH-1:0] c_out611;
output [32*C_WIDTH-1:0] c_out612;
output [32*C_WIDTH-1:0] c_out613;
output [32*C_WIDTH-1:0] c_out614;
output [32*C_WIDTH-1:0] c_out615;
output [32*C_WIDTH-1:0] c_out616;
output [32*C_WIDTH-1:0] c_out617;
output [32*C_WIDTH-1:0] c_out618;
output [32*C_WIDTH-1:0] c_out619;
output [32*C_WIDTH-1:0] c_out620;
output [32*C_WIDTH-1:0] c_out621;
output [32*C_WIDTH-1:0] c_out622;
output [32*C_WIDTH-1:0] c_out623;
output [32*C_WIDTH-1:0] c_out624;
output [32*C_WIDTH-1:0] c_out625;
output [32*C_WIDTH-1:0] c_out626;
output [32*C_WIDTH-1:0] c_out627;
output [32*C_WIDTH-1:0] c_out628;
output [32*C_WIDTH-1:0] c_out629;
output [32*C_WIDTH-1:0] c_out630;
output [32*C_WIDTH-1:0] c_out631;
output [32*C_WIDTH-1:0] c_out632;
output [32*C_WIDTH-1:0] c_out633;
output [32*C_WIDTH-1:0] c_out634;
output [32*C_WIDTH-1:0] c_out635;
output [32*C_WIDTH-1:0] c_out636;
output [32*C_WIDTH-1:0] c_out637;
output [32*C_WIDTH-1:0] c_out638;
output [32*C_WIDTH-1:0] c_out639;
output [32*C_WIDTH-1:0] c_out640;
output [32*C_WIDTH-1:0] c_out641;
output [32*C_WIDTH-1:0] c_out642;
output [32*C_WIDTH-1:0] c_out643;
output [32*C_WIDTH-1:0] c_out644;
output [32*C_WIDTH-1:0] c_out645;
output [32*C_WIDTH-1:0] c_out646;
output [32*C_WIDTH-1:0] c_out647;
output [32*C_WIDTH-1:0] c_out648;
output [32*C_WIDTH-1:0] c_out649;
output [32*C_WIDTH-1:0] c_out650;
output [32*C_WIDTH-1:0] c_out651;
output [32*C_WIDTH-1:0] c_out652;
output [32*C_WIDTH-1:0] c_out653;
output [32*C_WIDTH-1:0] c_out654;
output [32*C_WIDTH-1:0] c_out655;
output [32*C_WIDTH-1:0] c_out656;
output [32*C_WIDTH-1:0] c_out657;
output [32*C_WIDTH-1:0] c_out658;
output [32*C_WIDTH-1:0] c_out659;
output [32*C_WIDTH-1:0] c_out660;
output [32*C_WIDTH-1:0] c_out661;
output [32*C_WIDTH-1:0] c_out662;
output [32*C_WIDTH-1:0] c_out663;
output [32*C_WIDTH-1:0] c_out664;
output [32*C_WIDTH-1:0] c_out665;
output [32*C_WIDTH-1:0] c_out666;
output [32*C_WIDTH-1:0] c_out667;
output [32*C_WIDTH-1:0] c_out668;
output [32*C_WIDTH-1:0] c_out669;
output [32*C_WIDTH-1:0] c_out670;
output [32*C_WIDTH-1:0] c_out671;
output [32*C_WIDTH-1:0] c_out672;
output [32*C_WIDTH-1:0] c_out673;
output [32*C_WIDTH-1:0] c_out674;
output [32*C_WIDTH-1:0] c_out675;
output [32*C_WIDTH-1:0] c_out676;
output [32*C_WIDTH-1:0] c_out677;
output [32*C_WIDTH-1:0] c_out678;
output [32*C_WIDTH-1:0] c_out679;
output [32*C_WIDTH-1:0] c_out680;
output [32*C_WIDTH-1:0] c_out681;
output [32*C_WIDTH-1:0] c_out682;
output [32*C_WIDTH-1:0] c_out683;
output [32*C_WIDTH-1:0] c_out684;
output [32*C_WIDTH-1:0] c_out685;
output [32*C_WIDTH-1:0] c_out686;
output [32*C_WIDTH-1:0] c_out687;
output [32*C_WIDTH-1:0] c_out688;
output [32*C_WIDTH-1:0] c_out689;
output [32*C_WIDTH-1:0] c_out690;
output [32*C_WIDTH-1:0] c_out691;
output [32*C_WIDTH-1:0] c_out692;
output [32*C_WIDTH-1:0] c_out693;
output [32*C_WIDTH-1:0] c_out694;
output [32*C_WIDTH-1:0] c_out695;
output [32*C_WIDTH-1:0] c_out696;
output [32*C_WIDTH-1:0] c_out697;
output [32*C_WIDTH-1:0] c_out698;
output [32*C_WIDTH-1:0] c_out699;
output [32*C_WIDTH-1:0] c_out700;
output [32*C_WIDTH-1:0] c_out701;
output [32*C_WIDTH-1:0] c_out702;
output [32*C_WIDTH-1:0] c_out703;
output [32*C_WIDTH-1:0] c_out704;
output [32*C_WIDTH-1:0] c_out705;
output [32*C_WIDTH-1:0] c_out706;
output [32*C_WIDTH-1:0] c_out707;
output [32*C_WIDTH-1:0] c_out708;
output [32*C_WIDTH-1:0] c_out709;
output [32*C_WIDTH-1:0] c_out710;
output [32*C_WIDTH-1:0] c_out711;
output [32*C_WIDTH-1:0] c_out712;
output [32*C_WIDTH-1:0] c_out713;
output [32*C_WIDTH-1:0] c_out714;
output [32*C_WIDTH-1:0] c_out715;
output [32*C_WIDTH-1:0] c_out716;
output [32*C_WIDTH-1:0] c_out717;
output [32*C_WIDTH-1:0] c_out718;
output [32*C_WIDTH-1:0] c_out719;
output [32*C_WIDTH-1:0] c_out720;
output [32*C_WIDTH-1:0] c_out721;
output [32*C_WIDTH-1:0] c_out722;
output [32*C_WIDTH-1:0] c_out723;
output [32*C_WIDTH-1:0] c_out724;
output [32*C_WIDTH-1:0] c_out725;
output [32*C_WIDTH-1:0] c_out726;
output [32*C_WIDTH-1:0] c_out727;
output [32*C_WIDTH-1:0] c_out728;
output [32*C_WIDTH-1:0] c_out729;
output [32*C_WIDTH-1:0] c_out730;
output [32*C_WIDTH-1:0] c_out731;
output [32*C_WIDTH-1:0] c_out732;
output [32*C_WIDTH-1:0] c_out733;
output [32*C_WIDTH-1:0] c_out734;
output [32*C_WIDTH-1:0] c_out735;
output [32*C_WIDTH-1:0] c_out736;
output [32*C_WIDTH-1:0] c_out737;
output [32*C_WIDTH-1:0] c_out738;
output [32*C_WIDTH-1:0] c_out739;
output [32*C_WIDTH-1:0] c_out740;
output [32*C_WIDTH-1:0] c_out741;
output [32*C_WIDTH-1:0] c_out742;
output [32*C_WIDTH-1:0] c_out743;
output [32*C_WIDTH-1:0] c_out744;
output [32*C_WIDTH-1:0] c_out745;
output [32*C_WIDTH-1:0] c_out746;
output [32*C_WIDTH-1:0] c_out747;
output [32*C_WIDTH-1:0] c_out748;
output [32*C_WIDTH-1:0] c_out749;
output [32*C_WIDTH-1:0] c_out750;
output [32*C_WIDTH-1:0] c_out751;
output [32*C_WIDTH-1:0] c_out752;
output [32*C_WIDTH-1:0] c_out753;
output [32*C_WIDTH-1:0] c_out754;
output [32*C_WIDTH-1:0] c_out755;
output [32*C_WIDTH-1:0] c_out756;
output [32*C_WIDTH-1:0] c_out757;
output [32*C_WIDTH-1:0] c_out758;
output [32*C_WIDTH-1:0] c_out759;
output [32*C_WIDTH-1:0] c_out760;
output [32*C_WIDTH-1:0] c_out761;
output [32*C_WIDTH-1:0] c_out762;
output [32*C_WIDTH-1:0] c_out763;
output [32*C_WIDTH-1:0] c_out764;
output [32*C_WIDTH-1:0] c_out765;
output [32*C_WIDTH-1:0] c_out766;
output [32*C_WIDTH-1:0] c_out767;
output [32*C_WIDTH-1:0] c_out768;
output [32*C_WIDTH-1:0] c_out769;
output [32*C_WIDTH-1:0] c_out770;
output [32*C_WIDTH-1:0] c_out771;
output [32*C_WIDTH-1:0] c_out772;
output [32*C_WIDTH-1:0] c_out773;
output [32*C_WIDTH-1:0] c_out774;
output [32*C_WIDTH-1:0] c_out775;
output [32*C_WIDTH-1:0] c_out776;
output [32*C_WIDTH-1:0] c_out777;
output [32*C_WIDTH-1:0] c_out778;
output [32*C_WIDTH-1:0] c_out779;
output [32*C_WIDTH-1:0] c_out780;
output [32*C_WIDTH-1:0] c_out781;
output [32*C_WIDTH-1:0] c_out782;
output [32*C_WIDTH-1:0] c_out783;
output [32*C_WIDTH-1:0] c_out784;
output [32*C_WIDTH-1:0] c_out785;
output [32*C_WIDTH-1:0] c_out786;
output [32*C_WIDTH-1:0] c_out787;
output [32*C_WIDTH-1:0] c_out788;
output [32*C_WIDTH-1:0] c_out789;
output [32*C_WIDTH-1:0] c_out790;
output [32*C_WIDTH-1:0] c_out791;
output [32*C_WIDTH-1:0] c_out792;
output [32*C_WIDTH-1:0] c_out793;
output [32*C_WIDTH-1:0] c_out794;
output [32*C_WIDTH-1:0] c_out795;
output [32*C_WIDTH-1:0] c_out796;
output [32*C_WIDTH-1:0] c_out797;
output [32*C_WIDTH-1:0] c_out798;
output [32*C_WIDTH-1:0] c_out799;
output [32*C_WIDTH-1:0] c_out800;
output [32*C_WIDTH-1:0] c_out801;
output [32*C_WIDTH-1:0] c_out802;
output [32*C_WIDTH-1:0] c_out803;
output [32*C_WIDTH-1:0] c_out804;
output [32*C_WIDTH-1:0] c_out805;
output [32*C_WIDTH-1:0] c_out806;
output [32*C_WIDTH-1:0] c_out807;
output [32*C_WIDTH-1:0] c_out808;
output [32*C_WIDTH-1:0] c_out809;
output [32*C_WIDTH-1:0] c_out810;
output [32*C_WIDTH-1:0] c_out811;
output [32*C_WIDTH-1:0] c_out812;
output [32*C_WIDTH-1:0] c_out813;
output [32*C_WIDTH-1:0] c_out814;
output [32*C_WIDTH-1:0] c_out815;
output [32*C_WIDTH-1:0] c_out816;
output [32*C_WIDTH-1:0] c_out817;
output [32*C_WIDTH-1:0] c_out818;
output [32*C_WIDTH-1:0] c_out819;
output [32*C_WIDTH-1:0] c_out820;
output [32*C_WIDTH-1:0] c_out821;
output [32*C_WIDTH-1:0] c_out822;
output [32*C_WIDTH-1:0] c_out823;
output [32*C_WIDTH-1:0] c_out824;
output [32*C_WIDTH-1:0] c_out825;
output [32*C_WIDTH-1:0] c_out826;
output [32*C_WIDTH-1:0] c_out827;
output [32*C_WIDTH-1:0] c_out828;
output [32*C_WIDTH-1:0] c_out829;
output [32*C_WIDTH-1:0] c_out830;
output [32*C_WIDTH-1:0] c_out831;
output [32*C_WIDTH-1:0] c_out832;
output [32*C_WIDTH-1:0] c_out833;
output [32*C_WIDTH-1:0] c_out834;
output [32*C_WIDTH-1:0] c_out835;
output [32*C_WIDTH-1:0] c_out836;
output [32*C_WIDTH-1:0] c_out837;
output [32*C_WIDTH-1:0] c_out838;
output [32*C_WIDTH-1:0] c_out839;
output [32*C_WIDTH-1:0] c_out840;
output [32*C_WIDTH-1:0] c_out841;
output [32*C_WIDTH-1:0] c_out842;
output [32*C_WIDTH-1:0] c_out843;
output [32*C_WIDTH-1:0] c_out844;
output [32*C_WIDTH-1:0] c_out845;
output [32*C_WIDTH-1:0] c_out846;
output [32*C_WIDTH-1:0] c_out847;
output [32*C_WIDTH-1:0] c_out848;
output [32*C_WIDTH-1:0] c_out849;
output [32*C_WIDTH-1:0] c_out850;
output [32*C_WIDTH-1:0] c_out851;
output [32*C_WIDTH-1:0] c_out852;
output [32*C_WIDTH-1:0] c_out853;
output [32*C_WIDTH-1:0] c_out854;
output [32*C_WIDTH-1:0] c_out855;
output [32*C_WIDTH-1:0] c_out856;
output [32*C_WIDTH-1:0] c_out857;
output [32*C_WIDTH-1:0] c_out858;
output [32*C_WIDTH-1:0] c_out859;
output [32*C_WIDTH-1:0] c_out860;
output [32*C_WIDTH-1:0] c_out861;
output [32*C_WIDTH-1:0] c_out862;
output [32*C_WIDTH-1:0] c_out863;
output [32*C_WIDTH-1:0] c_out864;
output [32*C_WIDTH-1:0] c_out865;
output [32*C_WIDTH-1:0] c_out866;
output [32*C_WIDTH-1:0] c_out867;
output [32*C_WIDTH-1:0] c_out868;
output [32*C_WIDTH-1:0] c_out869;
output [32*C_WIDTH-1:0] c_out870;
output [32*C_WIDTH-1:0] c_out871;
output [32*C_WIDTH-1:0] c_out872;
output [32*C_WIDTH-1:0] c_out873;
output [32*C_WIDTH-1:0] c_out874;
output [32*C_WIDTH-1:0] c_out875;
output [32*C_WIDTH-1:0] c_out876;
output [32*C_WIDTH-1:0] c_out877;
output [32*C_WIDTH-1:0] c_out878;
output [32*C_WIDTH-1:0] c_out879;
output [32*C_WIDTH-1:0] c_out880;
output [32*C_WIDTH-1:0] c_out881;
output [32*C_WIDTH-1:0] c_out882;
output [32*C_WIDTH-1:0] c_out883;
output [32*C_WIDTH-1:0] c_out884;
output [32*C_WIDTH-1:0] c_out885;
output [32*C_WIDTH-1:0] c_out886;
output [32*C_WIDTH-1:0] c_out887;
output [32*C_WIDTH-1:0] c_out888;
output [32*C_WIDTH-1:0] c_out889;
output [32*C_WIDTH-1:0] c_out890;
output [32*C_WIDTH-1:0] c_out891;
output [32*C_WIDTH-1:0] c_out892;
output [32*C_WIDTH-1:0] c_out893;
output [32*C_WIDTH-1:0] c_out894;
output [32*C_WIDTH-1:0] c_out895;
output [32*C_WIDTH-1:0] c_out896;
output [32*C_WIDTH-1:0] c_out897;
output [32*C_WIDTH-1:0] c_out898;
output [32*C_WIDTH-1:0] c_out899;
output [32*C_WIDTH-1:0] c_out900;
output [32*C_WIDTH-1:0] c_out901;
output [32*C_WIDTH-1:0] c_out902;
output [32*C_WIDTH-1:0] c_out903;
output [32*C_WIDTH-1:0] c_out904;
output [32*C_WIDTH-1:0] c_out905;
output [32*C_WIDTH-1:0] c_out906;
output [32*C_WIDTH-1:0] c_out907;
output [32*C_WIDTH-1:0] c_out908;
output [32*C_WIDTH-1:0] c_out909;
output [32*C_WIDTH-1:0] c_out910;
output [32*C_WIDTH-1:0] c_out911;
output [32*C_WIDTH-1:0] c_out912;
output [32*C_WIDTH-1:0] c_out913;
output [32*C_WIDTH-1:0] c_out914;
output [32*C_WIDTH-1:0] c_out915;
output [32*C_WIDTH-1:0] c_out916;
output [32*C_WIDTH-1:0] c_out917;
output [32*C_WIDTH-1:0] c_out918;
output [32*C_WIDTH-1:0] c_out919;
output [32*C_WIDTH-1:0] c_out920;
output [32*C_WIDTH-1:0] c_out921;
output [32*C_WIDTH-1:0] c_out922;
output [32*C_WIDTH-1:0] c_out923;
output [32*C_WIDTH-1:0] c_out924;
output [32*C_WIDTH-1:0] c_out925;
output [32*C_WIDTH-1:0] c_out926;
output [32*C_WIDTH-1:0] c_out927;
output [32*C_WIDTH-1:0] c_out928;
output [32*C_WIDTH-1:0] c_out929;
output [32*C_WIDTH-1:0] c_out930;
output [32*C_WIDTH-1:0] c_out931;
output [32*C_WIDTH-1:0] c_out932;
output [32*C_WIDTH-1:0] c_out933;
output [32*C_WIDTH-1:0] c_out934;
output [32*C_WIDTH-1:0] c_out935;
output [32*C_WIDTH-1:0] c_out936;
output [32*C_WIDTH-1:0] c_out937;
output [32*C_WIDTH-1:0] c_out938;
output [32*C_WIDTH-1:0] c_out939;
output [32*C_WIDTH-1:0] c_out940;
output [32*C_WIDTH-1:0] c_out941;
output [32*C_WIDTH-1:0] c_out942;
output [32*C_WIDTH-1:0] c_out943;
output [32*C_WIDTH-1:0] c_out944;
output [32*C_WIDTH-1:0] c_out945;
output [32*C_WIDTH-1:0] c_out946;
output [32*C_WIDTH-1:0] c_out947;
output [32*C_WIDTH-1:0] c_out948;
output [32*C_WIDTH-1:0] c_out949;
output [32*C_WIDTH-1:0] c_out950;
output [32*C_WIDTH-1:0] c_out951;
output [32*C_WIDTH-1:0] c_out952;
output [32*C_WIDTH-1:0] c_out953;
output [32*C_WIDTH-1:0] c_out954;
output [32*C_WIDTH-1:0] c_out955;
output [32*C_WIDTH-1:0] c_out956;
output [32*C_WIDTH-1:0] c_out957;
output [32*C_WIDTH-1:0] c_out958;
output [32*C_WIDTH-1:0] c_out959;
output [32*C_WIDTH-1:0] c_out960;
output [32*C_WIDTH-1:0] c_out961;
output [32*C_WIDTH-1:0] c_out962;
output [32*C_WIDTH-1:0] c_out963;
output [32*C_WIDTH-1:0] c_out964;
output [32*C_WIDTH-1:0] c_out965;
output [32*C_WIDTH-1:0] c_out966;
output [32*C_WIDTH-1:0] c_out967;
output [32*C_WIDTH-1:0] c_out968;
output [32*C_WIDTH-1:0] c_out969;
output [32*C_WIDTH-1:0] c_out970;
output [32*C_WIDTH-1:0] c_out971;
output [32*C_WIDTH-1:0] c_out972;
output [32*C_WIDTH-1:0] c_out973;
output [32*C_WIDTH-1:0] c_out974;
output [32*C_WIDTH-1:0] c_out975;
output [32*C_WIDTH-1:0] c_out976;
output [32*C_WIDTH-1:0] c_out977;
output [32*C_WIDTH-1:0] c_out978;
output [32*C_WIDTH-1:0] c_out979;
output [32*C_WIDTH-1:0] c_out980;
output [32*C_WIDTH-1:0] c_out981;
output [32*C_WIDTH-1:0] c_out982;
output [32*C_WIDTH-1:0] c_out983;
output [32*C_WIDTH-1:0] c_out984;
output [32*C_WIDTH-1:0] c_out985;
output [32*C_WIDTH-1:0] c_out986;
output [32*C_WIDTH-1:0] c_out987;
output [32*C_WIDTH-1:0] c_out988;
output [32*C_WIDTH-1:0] c_out989;
output [32*C_WIDTH-1:0] c_out990;
output [32*C_WIDTH-1:0] c_out991;
output [32*C_WIDTH-1:0] c_out992;
output [32*C_WIDTH-1:0] c_out993;
output [32*C_WIDTH-1:0] c_out994;
output [32*C_WIDTH-1:0] c_out995;
output [32*C_WIDTH-1:0] c_out996;
output [32*C_WIDTH-1:0] c_out997;
output [32*C_WIDTH-1:0] c_out998;
output [32*C_WIDTH-1:0] c_out999;
output [32*C_WIDTH-1:0] c_out1000;
output [32*C_WIDTH-1:0] c_out1001;
output [32*C_WIDTH-1:0] c_out1002;
output [32*C_WIDTH-1:0] c_out1003;
output [32*C_WIDTH-1:0] c_out1004;
output [32*C_WIDTH-1:0] c_out1005;
output [32*C_WIDTH-1:0] c_out1006;
output [32*C_WIDTH-1:0] c_out1007;
output [32*C_WIDTH-1:0] c_out1008;
output [32*C_WIDTH-1:0] c_out1009;
output [32*C_WIDTH-1:0] c_out1010;
output [32*C_WIDTH-1:0] c_out1011;
output [32*C_WIDTH-1:0] c_out1012;
output [32*C_WIDTH-1:0] c_out1013;
output [32*C_WIDTH-1:0] c_out1014;
output [32*C_WIDTH-1:0] c_out1015;
output [32*C_WIDTH-1:0] c_out1016;
output [32*C_WIDTH-1:0] c_out1017;
output [32*C_WIDTH-1:0] c_out1018;
output [32*C_WIDTH-1:0] c_out1019;
output [32*C_WIDTH-1:0] c_out1020;
output [32*C_WIDTH-1:0] c_out1021;
output [32*C_WIDTH-1:0] c_out1022;
output [32*C_WIDTH-1:0] c_out1023;
output [32*C_WIDTH-1:0] c_out1024;
output [32*C_WIDTH-1:0] c_out1025;
output [32*C_WIDTH-1:0] c_out1026;
output [32*C_WIDTH-1:0] c_out1027;
output [32*C_WIDTH-1:0] c_out1028;
output [32*C_WIDTH-1:0] c_out1029;
output [32*C_WIDTH-1:0] c_out1030;
output [32*C_WIDTH-1:0] c_out1031;
output [32*C_WIDTH-1:0] c_out1032;
output [32*C_WIDTH-1:0] c_out1033;
output [32*C_WIDTH-1:0] c_out1034;
output [32*C_WIDTH-1:0] c_out1035;
output [32*C_WIDTH-1:0] c_out1036;
output [32*C_WIDTH-1:0] c_out1037;
output [32*C_WIDTH-1:0] c_out1038;
output [32*C_WIDTH-1:0] c_out1039;
output [32*C_WIDTH-1:0] c_out1040;
output [32*C_WIDTH-1:0] c_out1041;
output [32*C_WIDTH-1:0] c_out1042;
output [32*C_WIDTH-1:0] c_out1043;
output [32*C_WIDTH-1:0] c_out1044;
output [32*C_WIDTH-1:0] c_out1045;
output [32*C_WIDTH-1:0] c_out1046;
output [32*C_WIDTH-1:0] c_out1047;
output [32*C_WIDTH-1:0] c_out1048;
output [32*C_WIDTH-1:0] c_out1049;
output [32*C_WIDTH-1:0] c_out1050;
output [32*C_WIDTH-1:0] c_out1051;
output [32*C_WIDTH-1:0] c_out1052;
output [32*C_WIDTH-1:0] c_out1053;
output [32*C_WIDTH-1:0] c_out1054;
output [32*C_WIDTH-1:0] c_out1055;
output [32*C_WIDTH-1:0] c_out1056;
output [32*C_WIDTH-1:0] c_out1057;
output [32*C_WIDTH-1:0] c_out1058;
output [32*C_WIDTH-1:0] c_out1059;
output [32*C_WIDTH-1:0] c_out1060;
output [32*C_WIDTH-1:0] c_out1061;
output [32*C_WIDTH-1:0] c_out1062;
output [32*C_WIDTH-1:0] c_out1063;
output [32*C_WIDTH-1:0] c_out1064;
output [32*C_WIDTH-1:0] c_out1065;
output [32*C_WIDTH-1:0] c_out1066;
output [32*C_WIDTH-1:0] c_out1067;
output [32*C_WIDTH-1:0] c_out1068;
output [32*C_WIDTH-1:0] c_out1069;
output [32*C_WIDTH-1:0] c_out1070;
output [32*C_WIDTH-1:0] c_out1071;
output [32*C_WIDTH-1:0] c_out1072;
output [32*C_WIDTH-1:0] c_out1073;
output [32*C_WIDTH-1:0] c_out1074;
output [32*C_WIDTH-1:0] c_out1075;
output [32*C_WIDTH-1:0] c_out1076;
output [32*C_WIDTH-1:0] c_out1077;
output [32*C_WIDTH-1:0] c_out1078;
output [32*C_WIDTH-1:0] c_out1079;
output [32*C_WIDTH-1:0] c_out1080;
output [32*C_WIDTH-1:0] c_out1081;
output [32*C_WIDTH-1:0] c_out1082;
output [32*C_WIDTH-1:0] c_out1083;
output [32*C_WIDTH-1:0] c_out1084;
output [32*C_WIDTH-1:0] c_out1085;
output [32*C_WIDTH-1:0] c_out1086;
output [32*C_WIDTH-1:0] c_out1087;
output [32*C_WIDTH-1:0] c_out1088;
output [32*C_WIDTH-1:0] c_out1089;
output [32*C_WIDTH-1:0] c_out1090;
output [32*C_WIDTH-1:0] c_out1091;
output [32*C_WIDTH-1:0] c_out1092;
output [32*C_WIDTH-1:0] c_out1093;
output [32*C_WIDTH-1:0] c_out1094;
output [32*C_WIDTH-1:0] c_out1095;
output [32*C_WIDTH-1:0] c_out1096;
output [32*C_WIDTH-1:0] c_out1097;
output [32*C_WIDTH-1:0] c_out1098;
output [32*C_WIDTH-1:0] c_out1099;
output [32*C_WIDTH-1:0] c_out1100;
output [32*C_WIDTH-1:0] c_out1101;
output [32*C_WIDTH-1:0] c_out1102;
output [32*C_WIDTH-1:0] c_out1103;
output [32*C_WIDTH-1:0] c_out1104;
output [32*C_WIDTH-1:0] c_out1105;
output [32*C_WIDTH-1:0] c_out1106;
output [32*C_WIDTH-1:0] c_out1107;
output [32*C_WIDTH-1:0] c_out1108;
output [32*C_WIDTH-1:0] c_out1109;
output [32*C_WIDTH-1:0] c_out1110;
output [32*C_WIDTH-1:0] c_out1111;
output [32*C_WIDTH-1:0] c_out1112;
output [32*C_WIDTH-1:0] c_out1113;
output [32*C_WIDTH-1:0] c_out1114;
output [32*C_WIDTH-1:0] c_out1115;
output [32*C_WIDTH-1:0] c_out1116;
output [32*C_WIDTH-1:0] c_out1117;
output [32*C_WIDTH-1:0] c_out1118;
output [32*C_WIDTH-1:0] c_out1119;
output [32*C_WIDTH-1:0] c_out1120;
output [32*C_WIDTH-1:0] c_out1121;
output [32*C_WIDTH-1:0] c_out1122;
output [32*C_WIDTH-1:0] c_out1123;
output [32*C_WIDTH-1:0] c_out1124;
output [32*C_WIDTH-1:0] c_out1125;
output [32*C_WIDTH-1:0] c_out1126;
output [32*C_WIDTH-1:0] c_out1127;
output [32*C_WIDTH-1:0] c_out1128;
output [32*C_WIDTH-1:0] c_out1129;
output [32*C_WIDTH-1:0] c_out1130;
output [32*C_WIDTH-1:0] c_out1131;
output [32*C_WIDTH-1:0] c_out1132;
output [32*C_WIDTH-1:0] c_out1133;
output [32*C_WIDTH-1:0] c_out1134;
output [32*C_WIDTH-1:0] c_out1135;
output [32*C_WIDTH-1:0] c_out1136;
output [32*C_WIDTH-1:0] c_out1137;
output [32*C_WIDTH-1:0] c_out1138;
output [32*C_WIDTH-1:0] c_out1139;
output [32*C_WIDTH-1:0] c_out1140;
output [32*C_WIDTH-1:0] c_out1141;
output [32*C_WIDTH-1:0] c_out1142;
output [32*C_WIDTH-1:0] c_out1143;
output [32*C_WIDTH-1:0] c_out1144;
output [32*C_WIDTH-1:0] c_out1145;
output [32*C_WIDTH-1:0] c_out1146;
output [32*C_WIDTH-1:0] c_out1147;
output [32*C_WIDTH-1:0] c_out1148;
output [32*C_WIDTH-1:0] c_out1149;
output [32*C_WIDTH-1:0] c_out1150;
output [32*C_WIDTH-1:0] c_out1151;
output [32*C_WIDTH-1:0] c_out1152;
output [32*C_WIDTH-1:0] c_out1153;
output [32*C_WIDTH-1:0] c_out1154;
output [32*C_WIDTH-1:0] c_out1155;
output [32*C_WIDTH-1:0] c_out1156;
output [32*C_WIDTH-1:0] c_out1157;
output [32*C_WIDTH-1:0] c_out1158;
output [32*C_WIDTH-1:0] c_out1159;
output [32*C_WIDTH-1:0] c_out1160;
output [32*C_WIDTH-1:0] c_out1161;
output [32*C_WIDTH-1:0] c_out1162;
output [32*C_WIDTH-1:0] c_out1163;
output [32*C_WIDTH-1:0] c_out1164;
output [32*C_WIDTH-1:0] c_out1165;
output [32*C_WIDTH-1:0] c_out1166;
output [32*C_WIDTH-1:0] c_out1167;
output [32*C_WIDTH-1:0] c_out1168;
output [32*C_WIDTH-1:0] c_out1169;
output [32*C_WIDTH-1:0] c_out1170;
output [32*C_WIDTH-1:0] c_out1171;
output [32*C_WIDTH-1:0] c_out1172;
output [32*C_WIDTH-1:0] c_out1173;
output [32*C_WIDTH-1:0] c_out1174;
output [32*C_WIDTH-1:0] c_out1175;
output [32*C_WIDTH-1:0] c_out1176;
output [32*C_WIDTH-1:0] c_out1177;
output [32*C_WIDTH-1:0] c_out1178;
output [32*C_WIDTH-1:0] c_out1179;
output [32*C_WIDTH-1:0] c_out1180;
output [32*C_WIDTH-1:0] c_out1181;
output [32*C_WIDTH-1:0] c_out1182;
output [32*C_WIDTH-1:0] c_out1183;
output [32*C_WIDTH-1:0] c_out1184;
output [32*C_WIDTH-1:0] c_out1185;
output [32*C_WIDTH-1:0] c_out1186;
output [32*C_WIDTH-1:0] c_out1187;
output [32*C_WIDTH-1:0] c_out1188;
output [32*C_WIDTH-1:0] c_out1189;
output [32*C_WIDTH-1:0] c_out1190;
output [32*C_WIDTH-1:0] c_out1191;
output [32*C_WIDTH-1:0] c_out1192;
output [32*C_WIDTH-1:0] c_out1193;
output [32*C_WIDTH-1:0] c_out1194;
output [32*C_WIDTH-1:0] c_out1195;
output [32*C_WIDTH-1:0] c_out1196;
output [32*C_WIDTH-1:0] c_out1197;
output [32*C_WIDTH-1:0] c_out1198;
output [32*C_WIDTH-1:0] c_out1199;
output [32*C_WIDTH-1:0] c_out1200;
output [32*C_WIDTH-1:0] c_out1201;
output [32*C_WIDTH-1:0] c_out1202;
output [32*C_WIDTH-1:0] c_out1203;
output [32*C_WIDTH-1:0] c_out1204;
output [32*C_WIDTH-1:0] c_out1205;
output [32*C_WIDTH-1:0] c_out1206;
output [32*C_WIDTH-1:0] c_out1207;
output [32*C_WIDTH-1:0] c_out1208;
output [32*C_WIDTH-1:0] c_out1209;
output [32*C_WIDTH-1:0] c_out1210;
output [32*C_WIDTH-1:0] c_out1211;
output [32*C_WIDTH-1:0] c_out1212;
output [32*C_WIDTH-1:0] c_out1213;
output [32*C_WIDTH-1:0] c_out1214;
output [32*C_WIDTH-1:0] c_out1215;
output [32*C_WIDTH-1:0] c_out1216;
output [32*C_WIDTH-1:0] c_out1217;
output [32*C_WIDTH-1:0] c_out1218;
output [32*C_WIDTH-1:0] c_out1219;
output [32*C_WIDTH-1:0] c_out1220;
output [32*C_WIDTH-1:0] c_out1221;
output [32*C_WIDTH-1:0] c_out1222;
output [32*C_WIDTH-1:0] c_out1223;
output [32*C_WIDTH-1:0] c_out1224;
output [32*C_WIDTH-1:0] c_out1225;
output [32*C_WIDTH-1:0] c_out1226;
output [32*C_WIDTH-1:0] c_out1227;
output [32*C_WIDTH-1:0] c_out1228;
output [32*C_WIDTH-1:0] c_out1229;
output [32*C_WIDTH-1:0] c_out1230;
output [32*C_WIDTH-1:0] c_out1231;
output [32*C_WIDTH-1:0] c_out1232;
output [32*C_WIDTH-1:0] c_out1233;
output [32*C_WIDTH-1:0] c_out1234;
output [32*C_WIDTH-1:0] c_out1235;
output [32*C_WIDTH-1:0] c_out1236;
output [32*C_WIDTH-1:0] c_out1237;
output [32*C_WIDTH-1:0] c_out1238;
output [32*C_WIDTH-1:0] c_out1239;
output [32*C_WIDTH-1:0] c_out1240;
output [32*C_WIDTH-1:0] c_out1241;
output [32*C_WIDTH-1:0] c_out1242;
output [32*C_WIDTH-1:0] c_out1243;
output [32*C_WIDTH-1:0] c_out1244;
output [32*C_WIDTH-1:0] c_out1245;
output [32*C_WIDTH-1:0] c_out1246;
output [32*C_WIDTH-1:0] c_out1247;
output [32*C_WIDTH-1:0] c_out1248;
output [32*C_WIDTH-1:0] c_out1249;
output [32*C_WIDTH-1:0] c_out1250;
output [32*C_WIDTH-1:0] c_out1251;
output [32*C_WIDTH-1:0] c_out1252;
output [32*C_WIDTH-1:0] c_out1253;
output [32*C_WIDTH-1:0] c_out1254;
output [32*C_WIDTH-1:0] c_out1255;
output [32*C_WIDTH-1:0] c_out1256;
output [32*C_WIDTH-1:0] c_out1257;
output [32*C_WIDTH-1:0] c_out1258;
output [32*C_WIDTH-1:0] c_out1259;
output [32*C_WIDTH-1:0] c_out1260;
output [32*C_WIDTH-1:0] c_out1261;
output [32*C_WIDTH-1:0] c_out1262;
output [32*C_WIDTH-1:0] c_out1263;
output [32*C_WIDTH-1:0] c_out1264;
output [32*C_WIDTH-1:0] c_out1265;
output [32*C_WIDTH-1:0] c_out1266;
output [32*C_WIDTH-1:0] c_out1267;
output [32*C_WIDTH-1:0] c_out1268;
output [32*C_WIDTH-1:0] c_out1269;
output [32*C_WIDTH-1:0] c_out1270;
output [32*C_WIDTH-1:0] c_out1271;
output [32*C_WIDTH-1:0] c_out1272;
output [32*C_WIDTH-1:0] c_out1273;
output [32*C_WIDTH-1:0] c_out1274;
output [32*C_WIDTH-1:0] c_out1275;
output [32*C_WIDTH-1:0] c_out1276;
output [32*C_WIDTH-1:0] c_out1277;
output [32*C_WIDTH-1:0] c_out1278;
output [32*C_WIDTH-1:0] c_out1279;
output [32*C_WIDTH-1:0] c_out1280;
output [32*C_WIDTH-1:0] c_out1281;
output [32*C_WIDTH-1:0] c_out1282;
output [32*C_WIDTH-1:0] c_out1283;
output [32*C_WIDTH-1:0] c_out1284;
output [32*C_WIDTH-1:0] c_out1285;
output [32*C_WIDTH-1:0] c_out1286;
output [32*C_WIDTH-1:0] c_out1287;
output [32*C_WIDTH-1:0] c_out1288;
output [32*C_WIDTH-1:0] c_out1289;
output [32*C_WIDTH-1:0] c_out1290;
output [32*C_WIDTH-1:0] c_out1291;
output [32*C_WIDTH-1:0] c_out1292;
output [32*C_WIDTH-1:0] c_out1293;
output [32*C_WIDTH-1:0] c_out1294;
output [32*C_WIDTH-1:0] c_out1295;
output [32*C_WIDTH-1:0] c_out1296;
output [32*C_WIDTH-1:0] c_out1297;
output [32*C_WIDTH-1:0] c_out1298;
output [32*C_WIDTH-1:0] c_out1299;
output [32*C_WIDTH-1:0] c_out1300;
output [32*C_WIDTH-1:0] c_out1301;
output [32*C_WIDTH-1:0] c_out1302;
output [32*C_WIDTH-1:0] c_out1303;
output [32*C_WIDTH-1:0] c_out1304;
output [32*C_WIDTH-1:0] c_out1305;
output [32*C_WIDTH-1:0] c_out1306;
output [32*C_WIDTH-1:0] c_out1307;
output [32*C_WIDTH-1:0] c_out1308;
output [32*C_WIDTH-1:0] c_out1309;
output [32*C_WIDTH-1:0] c_out1310;
output [32*C_WIDTH-1:0] c_out1311;
output [32*C_WIDTH-1:0] c_out1312;
output [32*C_WIDTH-1:0] c_out1313;
output [32*C_WIDTH-1:0] c_out1314;
output [32*C_WIDTH-1:0] c_out1315;
output [32*C_WIDTH-1:0] c_out1316;
output [32*C_WIDTH-1:0] c_out1317;
output [32*C_WIDTH-1:0] c_out1318;
output [32*C_WIDTH-1:0] c_out1319;
output [32*C_WIDTH-1:0] c_out1320;
output [32*C_WIDTH-1:0] c_out1321;
output [32*C_WIDTH-1:0] c_out1322;
output [32*C_WIDTH-1:0] c_out1323;
output [32*C_WIDTH-1:0] c_out1324;
output [32*C_WIDTH-1:0] c_out1325;
output [32*C_WIDTH-1:0] c_out1326;
output [32*C_WIDTH-1:0] c_out1327;
output [32*C_WIDTH-1:0] c_out1328;
output [32*C_WIDTH-1:0] c_out1329;
output [32*C_WIDTH-1:0] c_out1330;
output [32*C_WIDTH-1:0] c_out1331;
output [32*C_WIDTH-1:0] c_out1332;
output [32*C_WIDTH-1:0] c_out1333;
output [32*C_WIDTH-1:0] c_out1334;
output [32*C_WIDTH-1:0] c_out1335;
output [32*C_WIDTH-1:0] c_out1336;
output [32*C_WIDTH-1:0] c_out1337;
output [32*C_WIDTH-1:0] c_out1338;
output [32*C_WIDTH-1:0] c_out1339;
output [32*C_WIDTH-1:0] c_out1340;
output [32*C_WIDTH-1:0] c_out1341;
output [32*C_WIDTH-1:0] c_out1342;
output [32*C_WIDTH-1:0] c_out1343;
output [32*C_WIDTH-1:0] c_out1344;
output [32*C_WIDTH-1:0] c_out1345;
output [32*C_WIDTH-1:0] c_out1346;
output [32*C_WIDTH-1:0] c_out1347;
output [32*C_WIDTH-1:0] c_out1348;
output [32*C_WIDTH-1:0] c_out1349;
output [32*C_WIDTH-1:0] c_out1350;
output [32*C_WIDTH-1:0] c_out1351;
output [32*C_WIDTH-1:0] c_out1352;
output [32*C_WIDTH-1:0] c_out1353;
output [32*C_WIDTH-1:0] c_out1354;
output [32*C_WIDTH-1:0] c_out1355;
output [32*C_WIDTH-1:0] c_out1356;
output [32*C_WIDTH-1:0] c_out1357;
output [32*C_WIDTH-1:0] c_out1358;
output [32*C_WIDTH-1:0] c_out1359;
output [32*C_WIDTH-1:0] c_out1360;
output [32*C_WIDTH-1:0] c_out1361;
output [32*C_WIDTH-1:0] c_out1362;
output [32*C_WIDTH-1:0] c_out1363;
output [32*C_WIDTH-1:0] c_out1364;
output [32*C_WIDTH-1:0] c_out1365;
output [32*C_WIDTH-1:0] c_out1366;
output [32*C_WIDTH-1:0] c_out1367;
output [32*C_WIDTH-1:0] c_out1368;
output [32*C_WIDTH-1:0] c_out1369;
output [32*C_WIDTH-1:0] c_out1370;
output [32*C_WIDTH-1:0] c_out1371;
output [32*C_WIDTH-1:0] c_out1372;
output [32*C_WIDTH-1:0] c_out1373;
output [32*C_WIDTH-1:0] c_out1374;
output [32*C_WIDTH-1:0] c_out1375;
output [32*C_WIDTH-1:0] c_out1376;
output [32*C_WIDTH-1:0] c_out1377;
output [32*C_WIDTH-1:0] c_out1378;
output [32*C_WIDTH-1:0] c_out1379;
output [32*C_WIDTH-1:0] c_out1380;
output [32*C_WIDTH-1:0] c_out1381;
output [32*C_WIDTH-1:0] c_out1382;
output [32*C_WIDTH-1:0] c_out1383;
output [32*C_WIDTH-1:0] c_out1384;
output [32*C_WIDTH-1:0] c_out1385;
output [32*C_WIDTH-1:0] c_out1386;
output [32*C_WIDTH-1:0] c_out1387;
output [32*C_WIDTH-1:0] c_out1388;
output [32*C_WIDTH-1:0] c_out1389;
output [32*C_WIDTH-1:0] c_out1390;
output [32*C_WIDTH-1:0] c_out1391;
output [32*C_WIDTH-1:0] c_out1392;
output [32*C_WIDTH-1:0] c_out1393;
output [32*C_WIDTH-1:0] c_out1394;
output [32*C_WIDTH-1:0] c_out1395;
output [32*C_WIDTH-1:0] c_out1396;
output [32*C_WIDTH-1:0] c_out1397;
output [32*C_WIDTH-1:0] c_out1398;
output [32*C_WIDTH-1:0] c_out1399;
output [32*C_WIDTH-1:0] c_out1400;
output [32*C_WIDTH-1:0] c_out1401;
output [32*C_WIDTH-1:0] c_out1402;
output [32*C_WIDTH-1:0] c_out1403;
output [32*C_WIDTH-1:0] c_out1404;
output [32*C_WIDTH-1:0] c_out1405;
output [32*C_WIDTH-1:0] c_out1406;
output [32*C_WIDTH-1:0] c_out1407;
output [32*C_WIDTH-1:0] c_out1408;
output [32*C_WIDTH-1:0] c_out1409;
output [32*C_WIDTH-1:0] c_out1410;
output [32*C_WIDTH-1:0] c_out1411;
output [32*C_WIDTH-1:0] c_out1412;
output [32*C_WIDTH-1:0] c_out1413;
output [32*C_WIDTH-1:0] c_out1414;
output [32*C_WIDTH-1:0] c_out1415;
output [32*C_WIDTH-1:0] c_out1416;
output [32*C_WIDTH-1:0] c_out1417;
output [32*C_WIDTH-1:0] c_out1418;
output [32*C_WIDTH-1:0] c_out1419;
output [32*C_WIDTH-1:0] c_out1420;
output [32*C_WIDTH-1:0] c_out1421;
output [32*C_WIDTH-1:0] c_out1422;
output [32*C_WIDTH-1:0] c_out1423;
output [32*C_WIDTH-1:0] c_out1424;
output [32*C_WIDTH-1:0] c_out1425;
output [32*C_WIDTH-1:0] c_out1426;
output [32*C_WIDTH-1:0] c_out1427;
output [32*C_WIDTH-1:0] c_out1428;
output [32*C_WIDTH-1:0] c_out1429;
output [32*C_WIDTH-1:0] c_out1430;
output [32*C_WIDTH-1:0] c_out1431;
output [32*C_WIDTH-1:0] c_out1432;
output [32*C_WIDTH-1:0] c_out1433;
output [32*C_WIDTH-1:0] c_out1434;
output [32*C_WIDTH-1:0] c_out1435;
output [32*C_WIDTH-1:0] c_out1436;
output [32*C_WIDTH-1:0] c_out1437;
output [32*C_WIDTH-1:0] c_out1438;
output [32*C_WIDTH-1:0] c_out1439;
output [32*C_WIDTH-1:0] c_out1440;
output [32*C_WIDTH-1:0] c_out1441;
output [32*C_WIDTH-1:0] c_out1442;
output [32*C_WIDTH-1:0] c_out1443;
output [32*C_WIDTH-1:0] c_out1444;
output [32*C_WIDTH-1:0] c_out1445;
output [32*C_WIDTH-1:0] c_out1446;
output [32*C_WIDTH-1:0] c_out1447;
output [32*C_WIDTH-1:0] c_out1448;
output [32*C_WIDTH-1:0] c_out1449;
output [32*C_WIDTH-1:0] c_out1450;
output [32*C_WIDTH-1:0] c_out1451;
output [32*C_WIDTH-1:0] c_out1452;
output [32*C_WIDTH-1:0] c_out1453;
output [32*C_WIDTH-1:0] c_out1454;
output [32*C_WIDTH-1:0] c_out1455;
output [32*C_WIDTH-1:0] c_out1456;
output [32*C_WIDTH-1:0] c_out1457;
output [32*C_WIDTH-1:0] c_out1458;
output [32*C_WIDTH-1:0] c_out1459;
output [32*C_WIDTH-1:0] c_out1460;
output [32*C_WIDTH-1:0] c_out1461;
output [32*C_WIDTH-1:0] c_out1462;
output [32*C_WIDTH-1:0] c_out1463;
output [32*C_WIDTH-1:0] c_out1464;
output [32*C_WIDTH-1:0] c_out1465;
output [32*C_WIDTH-1:0] c_out1466;
output [32*C_WIDTH-1:0] c_out1467;
output [32*C_WIDTH-1:0] c_out1468;
output [32*C_WIDTH-1:0] c_out1469;
output [32*C_WIDTH-1:0] c_out1470;
output [32*C_WIDTH-1:0] c_out1471;
output [32*C_WIDTH-1:0] c_out1472;
output [32*C_WIDTH-1:0] c_out1473;
output [32*C_WIDTH-1:0] c_out1474;
output [32*C_WIDTH-1:0] c_out1475;
output [32*C_WIDTH-1:0] c_out1476;
output [32*C_WIDTH-1:0] c_out1477;
output [32*C_WIDTH-1:0] c_out1478;
output [32*C_WIDTH-1:0] c_out1479;
output [32*C_WIDTH-1:0] c_out1480;
output [32*C_WIDTH-1:0] c_out1481;
output [32*C_WIDTH-1:0] c_out1482;
output [32*C_WIDTH-1:0] c_out1483;
output [32*C_WIDTH-1:0] c_out1484;
output [32*C_WIDTH-1:0] c_out1485;
output [32*C_WIDTH-1:0] c_out1486;
output [32*C_WIDTH-1:0] c_out1487;
output [32*C_WIDTH-1:0] c_out1488;
output [32*C_WIDTH-1:0] c_out1489;
output [32*C_WIDTH-1:0] c_out1490;
output [32*C_WIDTH-1:0] c_out1491;
output [32*C_WIDTH-1:0] c_out1492;
output [32*C_WIDTH-1:0] c_out1493;
output [32*C_WIDTH-1:0] c_out1494;
output [32*C_WIDTH-1:0] c_out1495;
output [32*C_WIDTH-1:0] c_out1496;
output [32*C_WIDTH-1:0] c_out1497;
output [32*C_WIDTH-1:0] c_out1498;
output [32*C_WIDTH-1:0] c_out1499;
output [32*C_WIDTH-1:0] c_out1500;
output [32*C_WIDTH-1:0] c_out1501;
output [32*C_WIDTH-1:0] c_out1502;
output [32*C_WIDTH-1:0] c_out1503;
output [32*C_WIDTH-1:0] c_out1504;
output [32*C_WIDTH-1:0] c_out1505;
output [32*C_WIDTH-1:0] c_out1506;
output [32*C_WIDTH-1:0] c_out1507;
output [32*C_WIDTH-1:0] c_out1508;
output [32*C_WIDTH-1:0] c_out1509;
output [32*C_WIDTH-1:0] c_out1510;
output [32*C_WIDTH-1:0] c_out1511;
output [32*C_WIDTH-1:0] c_out1512;
output [32*C_WIDTH-1:0] c_out1513;
output [32*C_WIDTH-1:0] c_out1514;
output [32*C_WIDTH-1:0] c_out1515;
output [32*C_WIDTH-1:0] c_out1516;
output [32*C_WIDTH-1:0] c_out1517;
output [32*C_WIDTH-1:0] c_out1518;
output [32*C_WIDTH-1:0] c_out1519;
output [32*C_WIDTH-1:0] c_out1520;
output [32*C_WIDTH-1:0] c_out1521;
output [32*C_WIDTH-1:0] c_out1522;
output [32*C_WIDTH-1:0] c_out1523;
output [32*C_WIDTH-1:0] c_out1524;
output [32*C_WIDTH-1:0] c_out1525;
output [32*C_WIDTH-1:0] c_out1526;
output [32*C_WIDTH-1:0] c_out1527;
output [32*C_WIDTH-1:0] c_out1528;
output [32*C_WIDTH-1:0] c_out1529;
output [32*C_WIDTH-1:0] c_out1530;
output [32*C_WIDTH-1:0] c_out1531;
output [32*C_WIDTH-1:0] c_out1532;
output [32*C_WIDTH-1:0] c_out1533;
output [32*C_WIDTH-1:0] c_out1534;
output [32*C_WIDTH-1:0] c_out1535;
output [32*C_WIDTH-1:0] c_out1536;
output [32*C_WIDTH-1:0] c_out1537;
output [32*C_WIDTH-1:0] c_out1538;
output [32*C_WIDTH-1:0] c_out1539;
output [32*C_WIDTH-1:0] c_out1540;
output [32*C_WIDTH-1:0] c_out1541;
output [32*C_WIDTH-1:0] c_out1542;
output [32*C_WIDTH-1:0] c_out1543;
output [32*C_WIDTH-1:0] c_out1544;
output [32*C_WIDTH-1:0] c_out1545;
output [32*C_WIDTH-1:0] c_out1546;
output [32*C_WIDTH-1:0] c_out1547;
output [32*C_WIDTH-1:0] c_out1548;
output [32*C_WIDTH-1:0] c_out1549;
output [32*C_WIDTH-1:0] c_out1550;
output [32*C_WIDTH-1:0] c_out1551;
output [32*C_WIDTH-1:0] c_out1552;
output [32*C_WIDTH-1:0] c_out1553;
output [32*C_WIDTH-1:0] c_out1554;
output [32*C_WIDTH-1:0] c_out1555;
output [32*C_WIDTH-1:0] c_out1556;
output [32*C_WIDTH-1:0] c_out1557;
output [32*C_WIDTH-1:0] c_out1558;
output [32*C_WIDTH-1:0] c_out1559;
output [32*C_WIDTH-1:0] c_out1560;
output [32*C_WIDTH-1:0] c_out1561;
output [32*C_WIDTH-1:0] c_out1562;
output [32*C_WIDTH-1:0] c_out1563;
output [32*C_WIDTH-1:0] c_out1564;
output [32*C_WIDTH-1:0] c_out1565;
output [32*C_WIDTH-1:0] c_out1566;
output [32*C_WIDTH-1:0] c_out1567;
output [32*C_WIDTH-1:0] c_out1568;
output [32*C_WIDTH-1:0] c_out1569;
output [32*C_WIDTH-1:0] c_out1570;
output [32*C_WIDTH-1:0] c_out1571;
output [32*C_WIDTH-1:0] c_out1572;
output [32*C_WIDTH-1:0] c_out1573;
output [32*C_WIDTH-1:0] c_out1574;
output [32*C_WIDTH-1:0] c_out1575;
output [32*C_WIDTH-1:0] c_out1576;
output [32*C_WIDTH-1:0] c_out1577;
output [32*C_WIDTH-1:0] c_out1578;
output [32*C_WIDTH-1:0] c_out1579;
output [32*C_WIDTH-1:0] c_out1580;
output [32*C_WIDTH-1:0] c_out1581;
output [32*C_WIDTH-1:0] c_out1582;
output [32*C_WIDTH-1:0] c_out1583;
output [32*C_WIDTH-1:0] c_out1584;
output [32*C_WIDTH-1:0] c_out1585;
output [32*C_WIDTH-1:0] c_out1586;
output [32*C_WIDTH-1:0] c_out1587;
output [32*C_WIDTH-1:0] c_out1588;
output [32*C_WIDTH-1:0] c_out1589;
output [32*C_WIDTH-1:0] c_out1590;
output [32*C_WIDTH-1:0] c_out1591;
output [32*C_WIDTH-1:0] c_out1592;
output [32*C_WIDTH-1:0] c_out1593;
output [32*C_WIDTH-1:0] c_out1594;
output [32*C_WIDTH-1:0] c_out1595;
output [32*C_WIDTH-1:0] c_out1596;
output [32*C_WIDTH-1:0] c_out1597;
output [32*C_WIDTH-1:0] c_out1598;
output [32*C_WIDTH-1:0] c_out1599;
output [32*C_WIDTH-1:0] c_out1600;
output [32*C_WIDTH-1:0] c_out1601;
output [32*C_WIDTH-1:0] c_out1602;
output [32*C_WIDTH-1:0] c_out1603;
output [32*C_WIDTH-1:0] c_out1604;
output [32*C_WIDTH-1:0] c_out1605;
output [32*C_WIDTH-1:0] c_out1606;
output [32*C_WIDTH-1:0] c_out1607;
output [32*C_WIDTH-1:0] c_out1608;
output [32*C_WIDTH-1:0] c_out1609;
output [32*C_WIDTH-1:0] c_out1610;
output [32*C_WIDTH-1:0] c_out1611;
output [32*C_WIDTH-1:0] c_out1612;
output [32*C_WIDTH-1:0] c_out1613;
output [32*C_WIDTH-1:0] c_out1614;
output [32*C_WIDTH-1:0] c_out1615;
output [32*C_WIDTH-1:0] c_out1616;
output [32*C_WIDTH-1:0] c_out1617;
output [32*C_WIDTH-1:0] c_out1618;
output [32*C_WIDTH-1:0] c_out1619;
output [32*C_WIDTH-1:0] c_out1620;
output [32*C_WIDTH-1:0] c_out1621;
output [32*C_WIDTH-1:0] c_out1622;
output [32*C_WIDTH-1:0] c_out1623;
output [32*C_WIDTH-1:0] c_out1624;
output [32*C_WIDTH-1:0] c_out1625;
output [32*C_WIDTH-1:0] c_out1626;
output [32*C_WIDTH-1:0] c_out1627;
output [32*C_WIDTH-1:0] c_out1628;
output [32*C_WIDTH-1:0] c_out1629;
output [32*C_WIDTH-1:0] c_out1630;
output [32*C_WIDTH-1:0] c_out1631;
output [32*C_WIDTH-1:0] c_out1632;
output [32*C_WIDTH-1:0] c_out1633;
output [32*C_WIDTH-1:0] c_out1634;
output [32*C_WIDTH-1:0] c_out1635;
output [32*C_WIDTH-1:0] c_out1636;
output [32*C_WIDTH-1:0] c_out1637;
output [32*C_WIDTH-1:0] c_out1638;
output [32*C_WIDTH-1:0] c_out1639;
output [32*C_WIDTH-1:0] c_out1640;
output [32*C_WIDTH-1:0] c_out1641;
output [32*C_WIDTH-1:0] c_out1642;
output [32*C_WIDTH-1:0] c_out1643;
output [32*C_WIDTH-1:0] c_out1644;
output [32*C_WIDTH-1:0] c_out1645;
output [32*C_WIDTH-1:0] c_out1646;
output [32*C_WIDTH-1:0] c_out1647;
output [32*C_WIDTH-1:0] c_out1648;
output [32*C_WIDTH-1:0] c_out1649;
output [32*C_WIDTH-1:0] c_out1650;
output [32*C_WIDTH-1:0] c_out1651;
output [32*C_WIDTH-1:0] c_out1652;
output [32*C_WIDTH-1:0] c_out1653;
output [32*C_WIDTH-1:0] c_out1654;
output [32*C_WIDTH-1:0] c_out1655;
output [32*C_WIDTH-1:0] c_out1656;
output [32*C_WIDTH-1:0] c_out1657;
output [32*C_WIDTH-1:0] c_out1658;
output [32*C_WIDTH-1:0] c_out1659;
output [32*C_WIDTH-1:0] c_out1660;
output [32*C_WIDTH-1:0] c_out1661;
output [32*C_WIDTH-1:0] c_out1662;
output [32*C_WIDTH-1:0] c_out1663;
output [32*C_WIDTH-1:0] c_out1664;
output [32*C_WIDTH-1:0] c_out1665;
output [32*C_WIDTH-1:0] c_out1666;
output [32*C_WIDTH-1:0] c_out1667;
output [32*C_WIDTH-1:0] c_out1668;
output [32*C_WIDTH-1:0] c_out1669;
output [32*C_WIDTH-1:0] c_out1670;
output [32*C_WIDTH-1:0] c_out1671;
output [32*C_WIDTH-1:0] c_out1672;
output [32*C_WIDTH-1:0] c_out1673;
output [32*C_WIDTH-1:0] c_out1674;
output [32*C_WIDTH-1:0] c_out1675;
output [32*C_WIDTH-1:0] c_out1676;
output [32*C_WIDTH-1:0] c_out1677;
output [32*C_WIDTH-1:0] c_out1678;
output [32*C_WIDTH-1:0] c_out1679;
output [32*C_WIDTH-1:0] c_out1680;
output [32*C_WIDTH-1:0] c_out1681;
output [32*C_WIDTH-1:0] c_out1682;
output [32*C_WIDTH-1:0] c_out1683;
output [32*C_WIDTH-1:0] c_out1684;
output [32*C_WIDTH-1:0] c_out1685;
output [32*C_WIDTH-1:0] c_out1686;
output [32*C_WIDTH-1:0] c_out1687;
output [32*C_WIDTH-1:0] c_out1688;
output [32*C_WIDTH-1:0] c_out1689;
output [32*C_WIDTH-1:0] c_out1690;
output [32*C_WIDTH-1:0] c_out1691;
output [32*C_WIDTH-1:0] c_out1692;
output [32*C_WIDTH-1:0] c_out1693;
output [32*C_WIDTH-1:0] c_out1694;
output [32*C_WIDTH-1:0] c_out1695;
output [32*C_WIDTH-1:0] c_out1696;
output [32*C_WIDTH-1:0] c_out1697;
output [32*C_WIDTH-1:0] c_out1698;
output [32*C_WIDTH-1:0] c_out1699;
output [32*C_WIDTH-1:0] c_out1700;
output [32*C_WIDTH-1:0] c_out1701;
output [32*C_WIDTH-1:0] c_out1702;
output [32*C_WIDTH-1:0] c_out1703;
output [32*C_WIDTH-1:0] c_out1704;
output [32*C_WIDTH-1:0] c_out1705;
output [32*C_WIDTH-1:0] c_out1706;
output [32*C_WIDTH-1:0] c_out1707;
output [32*C_WIDTH-1:0] c_out1708;
output [32*C_WIDTH-1:0] c_out1709;
output [32*C_WIDTH-1:0] c_out1710;
output [32*C_WIDTH-1:0] c_out1711;
output [32*C_WIDTH-1:0] c_out1712;
output [32*C_WIDTH-1:0] c_out1713;
output [32*C_WIDTH-1:0] c_out1714;
output [32*C_WIDTH-1:0] c_out1715;
output [32*C_WIDTH-1:0] c_out1716;
output [32*C_WIDTH-1:0] c_out1717;
output [32*C_WIDTH-1:0] c_out1718;
output [32*C_WIDTH-1:0] c_out1719;
output [32*C_WIDTH-1:0] c_out1720;
output [32*C_WIDTH-1:0] c_out1721;
output [32*C_WIDTH-1:0] c_out1722;
output [32*C_WIDTH-1:0] c_out1723;
output [32*C_WIDTH-1:0] c_out1724;
output [32*C_WIDTH-1:0] c_out1725;
output [32*C_WIDTH-1:0] c_out1726;
output [32*C_WIDTH-1:0] c_out1727;
output [32*C_WIDTH-1:0] c_out1728;
output [32*C_WIDTH-1:0] c_out1729;
output [32*C_WIDTH-1:0] c_out1730;
output [32*C_WIDTH-1:0] c_out1731;
output [32*C_WIDTH-1:0] c_out1732;
output [32*C_WIDTH-1:0] c_out1733;
output [32*C_WIDTH-1:0] c_out1734;
output [32*C_WIDTH-1:0] c_out1735;
output [32*C_WIDTH-1:0] c_out1736;
output [32*C_WIDTH-1:0] c_out1737;
output [32*C_WIDTH-1:0] c_out1738;
output [32*C_WIDTH-1:0] c_out1739;
output [32*C_WIDTH-1:0] c_out1740;
output [32*C_WIDTH-1:0] c_out1741;
output [32*C_WIDTH-1:0] c_out1742;
output [32*C_WIDTH-1:0] c_out1743;
output [32*C_WIDTH-1:0] c_out1744;
output [32*C_WIDTH-1:0] c_out1745;
output [32*C_WIDTH-1:0] c_out1746;
output [32*C_WIDTH-1:0] c_out1747;
output [32*C_WIDTH-1:0] c_out1748;
output [32*C_WIDTH-1:0] c_out1749;
output [32*C_WIDTH-1:0] c_out1750;
output [32*C_WIDTH-1:0] c_out1751;
output [32*C_WIDTH-1:0] c_out1752;
output [32*C_WIDTH-1:0] c_out1753;
output [32*C_WIDTH-1:0] c_out1754;
output [32*C_WIDTH-1:0] c_out1755;
output [32*C_WIDTH-1:0] c_out1756;
output [32*C_WIDTH-1:0] c_out1757;
output [32*C_WIDTH-1:0] c_out1758;
output [32*C_WIDTH-1:0] c_out1759;
output [32*C_WIDTH-1:0] c_out1760;
output [32*C_WIDTH-1:0] c_out1761;
output [32*C_WIDTH-1:0] c_out1762;
output [32*C_WIDTH-1:0] c_out1763;
output [32*C_WIDTH-1:0] c_out1764;
output [32*C_WIDTH-1:0] c_out1765;
output [32*C_WIDTH-1:0] c_out1766;
output [32*C_WIDTH-1:0] c_out1767;
output [32*C_WIDTH-1:0] c_out1768;
output [32*C_WIDTH-1:0] c_out1769;
output [32*C_WIDTH-1:0] c_out1770;
output [32*C_WIDTH-1:0] c_out1771;
output [32*C_WIDTH-1:0] c_out1772;
output [32*C_WIDTH-1:0] c_out1773;
output [32*C_WIDTH-1:0] c_out1774;
output [32*C_WIDTH-1:0] c_out1775;
output [32*C_WIDTH-1:0] c_out1776;
output [32*C_WIDTH-1:0] c_out1777;
output [32*C_WIDTH-1:0] c_out1778;
output [32*C_WIDTH-1:0] c_out1779;
output [32*C_WIDTH-1:0] c_out1780;
output [32*C_WIDTH-1:0] c_out1781;
output [32*C_WIDTH-1:0] c_out1782;
output [32*C_WIDTH-1:0] c_out1783;
output [32*C_WIDTH-1:0] c_out1784;
output [32*C_WIDTH-1:0] c_out1785;
output [32*C_WIDTH-1:0] c_out1786;
output [32*C_WIDTH-1:0] c_out1787;
output [32*C_WIDTH-1:0] c_out1788;
output [32*C_WIDTH-1:0] c_out1789;
output [32*C_WIDTH-1:0] c_out1790;
output [32*C_WIDTH-1:0] c_out1791;
output [32*C_WIDTH-1:0] c_out1792;
output [32*C_WIDTH-1:0] c_out1793;
output [32*C_WIDTH-1:0] c_out1794;
output [32*C_WIDTH-1:0] c_out1795;
output [32*C_WIDTH-1:0] c_out1796;
output [32*C_WIDTH-1:0] c_out1797;
output [32*C_WIDTH-1:0] c_out1798;
output [32*C_WIDTH-1:0] c_out1799;
output [32*C_WIDTH-1:0] c_out1800;
output [32*C_WIDTH-1:0] c_out1801;
output [32*C_WIDTH-1:0] c_out1802;
output [32*C_WIDTH-1:0] c_out1803;
output [32*C_WIDTH-1:0] c_out1804;
output [32*C_WIDTH-1:0] c_out1805;
output [32*C_WIDTH-1:0] c_out1806;
output [32*C_WIDTH-1:0] c_out1807;
output [32*C_WIDTH-1:0] c_out1808;
output [32*C_WIDTH-1:0] c_out1809;
output [32*C_WIDTH-1:0] c_out1810;
output [32*C_WIDTH-1:0] c_out1811;
output [32*C_WIDTH-1:0] c_out1812;
output [32*C_WIDTH-1:0] c_out1813;
output [32*C_WIDTH-1:0] c_out1814;
output [32*C_WIDTH-1:0] c_out1815;
output [32*C_WIDTH-1:0] c_out1816;
output [32*C_WIDTH-1:0] c_out1817;
output [32*C_WIDTH-1:0] c_out1818;
output [32*C_WIDTH-1:0] c_out1819;
output [32*C_WIDTH-1:0] c_out1820;
output [32*C_WIDTH-1:0] c_out1821;
output [32*C_WIDTH-1:0] c_out1822;
output [32*C_WIDTH-1:0] c_out1823;
output [32*C_WIDTH-1:0] c_out1824;
output [32*C_WIDTH-1:0] c_out1825;
output [32*C_WIDTH-1:0] c_out1826;
output [32*C_WIDTH-1:0] c_out1827;
output [32*C_WIDTH-1:0] c_out1828;
output [32*C_WIDTH-1:0] c_out1829;
output [32*C_WIDTH-1:0] c_out1830;
output [32*C_WIDTH-1:0] c_out1831;
output [32*C_WIDTH-1:0] c_out1832;
output [32*C_WIDTH-1:0] c_out1833;
output [32*C_WIDTH-1:0] c_out1834;
output [32*C_WIDTH-1:0] c_out1835;
output [32*C_WIDTH-1:0] c_out1836;
output [32*C_WIDTH-1:0] c_out1837;
output [32*C_WIDTH-1:0] c_out1838;
output [32*C_WIDTH-1:0] c_out1839;
output [32*C_WIDTH-1:0] c_out1840;
output [32*C_WIDTH-1:0] c_out1841;
output [32*C_WIDTH-1:0] c_out1842;
output [32*C_WIDTH-1:0] c_out1843;
output [32*C_WIDTH-1:0] c_out1844;
output [32*C_WIDTH-1:0] c_out1845;
output [32*C_WIDTH-1:0] c_out1846;
output [32*C_WIDTH-1:0] c_out1847;
output [32*C_WIDTH-1:0] c_out1848;
output [32*C_WIDTH-1:0] c_out1849;
output [32*C_WIDTH-1:0] c_out1850;
output [32*C_WIDTH-1:0] c_out1851;
output [32*C_WIDTH-1:0] c_out1852;
output [32*C_WIDTH-1:0] c_out1853;
output [32*C_WIDTH-1:0] c_out1854;
output [32*C_WIDTH-1:0] c_out1855;
output [32*C_WIDTH-1:0] c_out1856;
output [32*C_WIDTH-1:0] c_out1857;
output [32*C_WIDTH-1:0] c_out1858;
output [32*C_WIDTH-1:0] c_out1859;
output [32*C_WIDTH-1:0] c_out1860;
output [32*C_WIDTH-1:0] c_out1861;
output [32*C_WIDTH-1:0] c_out1862;
output [32*C_WIDTH-1:0] c_out1863;
output [32*C_WIDTH-1:0] c_out1864;
output [32*C_WIDTH-1:0] c_out1865;
output [32*C_WIDTH-1:0] c_out1866;
output [32*C_WIDTH-1:0] c_out1867;
output [32*C_WIDTH-1:0] c_out1868;
output [32*C_WIDTH-1:0] c_out1869;
output [32*C_WIDTH-1:0] c_out1870;
output [32*C_WIDTH-1:0] c_out1871;
output [32*C_WIDTH-1:0] c_out1872;
output [32*C_WIDTH-1:0] c_out1873;
output [32*C_WIDTH-1:0] c_out1874;
output [32*C_WIDTH-1:0] c_out1875;
output [32*C_WIDTH-1:0] c_out1876;
output [32*C_WIDTH-1:0] c_out1877;
output [32*C_WIDTH-1:0] c_out1878;
output [32*C_WIDTH-1:0] c_out1879;
output [32*C_WIDTH-1:0] c_out1880;
output [32*C_WIDTH-1:0] c_out1881;
output [32*C_WIDTH-1:0] c_out1882;
output [32*C_WIDTH-1:0] c_out1883;
output [32*C_WIDTH-1:0] c_out1884;
output [32*C_WIDTH-1:0] c_out1885;
output [32*C_WIDTH-1:0] c_out1886;
output [32*C_WIDTH-1:0] c_out1887;
output [32*C_WIDTH-1:0] c_out1888;
output [32*C_WIDTH-1:0] c_out1889;
output [32*C_WIDTH-1:0] c_out1890;
output [32*C_WIDTH-1:0] c_out1891;
output [32*C_WIDTH-1:0] c_out1892;
output [32*C_WIDTH-1:0] c_out1893;
output [32*C_WIDTH-1:0] c_out1894;
output [32*C_WIDTH-1:0] c_out1895;
output [32*C_WIDTH-1:0] c_out1896;
output [32*C_WIDTH-1:0] c_out1897;
output [32*C_WIDTH-1:0] c_out1898;
output [32*C_WIDTH-1:0] c_out1899;
output [32*C_WIDTH-1:0] c_out1900;
output [32*C_WIDTH-1:0] c_out1901;
output [32*C_WIDTH-1:0] c_out1902;
output [32*C_WIDTH-1:0] c_out1903;
output [32*C_WIDTH-1:0] c_out1904;
output [32*C_WIDTH-1:0] c_out1905;
output [32*C_WIDTH-1:0] c_out1906;
output [32*C_WIDTH-1:0] c_out1907;
output [32*C_WIDTH-1:0] c_out1908;
output [32*C_WIDTH-1:0] c_out1909;
output [32*C_WIDTH-1:0] c_out1910;
output [32*C_WIDTH-1:0] c_out1911;
output [32*C_WIDTH-1:0] c_out1912;
output [32*C_WIDTH-1:0] c_out1913;
output [32*C_WIDTH-1:0] c_out1914;
output [32*C_WIDTH-1:0] c_out1915;
output [32*C_WIDTH-1:0] c_out1916;
output [32*C_WIDTH-1:0] c_out1917;
output [32*C_WIDTH-1:0] c_out1918;
output [32*C_WIDTH-1:0] c_out1919;
output [32*C_WIDTH-1:0] c_out1920;
output [32*C_WIDTH-1:0] c_out1921;
output [32*C_WIDTH-1:0] c_out1922;
output [32*C_WIDTH-1:0] c_out1923;
output [32*C_WIDTH-1:0] c_out1924;
output [32*C_WIDTH-1:0] c_out1925;
output [32*C_WIDTH-1:0] c_out1926;
output [32*C_WIDTH-1:0] c_out1927;
output [32*C_WIDTH-1:0] c_out1928;
output [32*C_WIDTH-1:0] c_out1929;
output [32*C_WIDTH-1:0] c_out1930;
output [32*C_WIDTH-1:0] c_out1931;
output [32*C_WIDTH-1:0] c_out1932;
output [32*C_WIDTH-1:0] c_out1933;
output [32*C_WIDTH-1:0] c_out1934;
output [32*C_WIDTH-1:0] c_out1935;
output [32*C_WIDTH-1:0] c_out1936;
output [32*C_WIDTH-1:0] c_out1937;
output [32*C_WIDTH-1:0] c_out1938;
output [32*C_WIDTH-1:0] c_out1939;
output [32*C_WIDTH-1:0] c_out1940;
output [32*C_WIDTH-1:0] c_out1941;
output [32*C_WIDTH-1:0] c_out1942;
output [32*C_WIDTH-1:0] c_out1943;
output [32*C_WIDTH-1:0] c_out1944;
output [32*C_WIDTH-1:0] c_out1945;
output [32*C_WIDTH-1:0] c_out1946;
output [32*C_WIDTH-1:0] c_out1947;
output [32*C_WIDTH-1:0] c_out1948;
output [32*C_WIDTH-1:0] c_out1949;
output [32*C_WIDTH-1:0] c_out1950;
output [32*C_WIDTH-1:0] c_out1951;
output [32*C_WIDTH-1:0] c_out1952;
output [32*C_WIDTH-1:0] c_out1953;
output [32*C_WIDTH-1:0] c_out1954;
output [32*C_WIDTH-1:0] c_out1955;
output [32*C_WIDTH-1:0] c_out1956;
output [32*C_WIDTH-1:0] c_out1957;
output [32*C_WIDTH-1:0] c_out1958;
output [32*C_WIDTH-1:0] c_out1959;
output [32*C_WIDTH-1:0] c_out1960;
output [32*C_WIDTH-1:0] c_out1961;
output [32*C_WIDTH-1:0] c_out1962;
output [32*C_WIDTH-1:0] c_out1963;
output [32*C_WIDTH-1:0] c_out1964;
output [32*C_WIDTH-1:0] c_out1965;
output [32*C_WIDTH-1:0] c_out1966;
output [32*C_WIDTH-1:0] c_out1967;
output [32*C_WIDTH-1:0] c_out1968;
output [32*C_WIDTH-1:0] c_out1969;
output [32*C_WIDTH-1:0] c_out1970;
output [32*C_WIDTH-1:0] c_out1971;
output [32*C_WIDTH-1:0] c_out1972;
output [32*C_WIDTH-1:0] c_out1973;
output [32*C_WIDTH-1:0] c_out1974;
output [32*C_WIDTH-1:0] c_out1975;
output [32*C_WIDTH-1:0] c_out1976;
output [32*C_WIDTH-1:0] c_out1977;
output [32*C_WIDTH-1:0] c_out1978;
output [32*C_WIDTH-1:0] c_out1979;
output [32*C_WIDTH-1:0] c_out1980;
output [32*C_WIDTH-1:0] c_out1981;
output [32*C_WIDTH-1:0] c_out1982;
output [32*C_WIDTH-1:0] c_out1983;
output [32*C_WIDTH-1:0] c_out1984;
output [32*C_WIDTH-1:0] c_out1985;
output [32*C_WIDTH-1:0] c_out1986;
output [32*C_WIDTH-1:0] c_out1987;
output [32*C_WIDTH-1:0] c_out1988;
output [32*C_WIDTH-1:0] c_out1989;
output [32*C_WIDTH-1:0] c_out1990;
output [32*C_WIDTH-1:0] c_out1991;
output [32*C_WIDTH-1:0] c_out1992;
output [32*C_WIDTH-1:0] c_out1993;
output [32*C_WIDTH-1:0] c_out1994;
output [32*C_WIDTH-1:0] c_out1995;
output [32*C_WIDTH-1:0] c_out1996;
output [32*C_WIDTH-1:0] c_out1997;
output [32*C_WIDTH-1:0] c_out1998;
output [32*C_WIDTH-1:0] c_out1999;
output [32*C_WIDTH-1:0] c_out2000;
output [32*C_WIDTH-1:0] c_out2001;
output [32*C_WIDTH-1:0] c_out2002;
output [32*C_WIDTH-1:0] c_out2003;
output [32*C_WIDTH-1:0] c_out2004;
output [32*C_WIDTH-1:0] c_out2005;
output [32*C_WIDTH-1:0] c_out2006;
output [32*C_WIDTH-1:0] c_out2007;
output [32*C_WIDTH-1:0] c_out2008;
output [32*C_WIDTH-1:0] c_out2009;
output [32*C_WIDTH-1:0] c_out2010;
output [32*C_WIDTH-1:0] c_out2011;
output [32*C_WIDTH-1:0] c_out2012;
output [32*C_WIDTH-1:0] c_out2013;
output [32*C_WIDTH-1:0] c_out2014;
output [32*C_WIDTH-1:0] c_out2015;
output [32*C_WIDTH-1:0] c_out2016;
output [32*C_WIDTH-1:0] c_out2017;
output [32*C_WIDTH-1:0] c_out2018;
output [32*C_WIDTH-1:0] c_out2019;
output [32*C_WIDTH-1:0] c_out2020;
output [32*C_WIDTH-1:0] c_out2021;
output [32*C_WIDTH-1:0] c_out2022;
output [32*C_WIDTH-1:0] c_out2023;
output [32*C_WIDTH-1:0] c_out2024;
output [32*C_WIDTH-1:0] c_out2025;
output [32*C_WIDTH-1:0] c_out2026;
output [32*C_WIDTH-1:0] c_out2027;
output [32*C_WIDTH-1:0] c_out2028;
output [32*C_WIDTH-1:0] c_out2029;
output [32*C_WIDTH-1:0] c_out2030;
output [32*C_WIDTH-1:0] c_out2031;
output [32*C_WIDTH-1:0] c_out2032;
output [32*C_WIDTH-1:0] c_out2033;
output [32*C_WIDTH-1:0] c_out2034;
output [32*C_WIDTH-1:0] c_out2035;
output [32*C_WIDTH-1:0] c_out2036;
output [32*C_WIDTH-1:0] c_out2037;
output [32*C_WIDTH-1:0] c_out2038;
output [32*C_WIDTH-1:0] c_out2039;
output [32*C_WIDTH-1:0] c_out2040;
output [32*C_WIDTH-1:0] c_out2041;
output [32*C_WIDTH-1:0] c_out2042;
output [32*C_WIDTH-1:0] c_out2043;
output [32*C_WIDTH-1:0] c_out2044;
output [32*C_WIDTH-1:0] c_out2045;
output [32*C_WIDTH-1:0] c_out2046;
output [32*C_WIDTH-1:0] c_out2047;
​

output [256*WIDTH-1:0] out_act;
output [256*WIDTH-1:0] out_weight;


wire [128*WIDTH-1:0] act_0;
wire [128*WIDTH-1:0] act_1;
wire [128*WIDTH-1:0] weight_0;
wire [128*WIDTH-1:0] weight_1;

wire [128*WIDTH-1:0] outact_0;
wire [128*WIDTH-1:0] outact_1;
wire [128*WIDTH-1:0] outweight_0;
wire [128*WIDTH-1:0] outweight_1;

wire [128*WIDTH-1:0] act0_1;
wire [128*WIDTH-1:0] act2_3;
wire [128*WIDTH-1:0] weight0_2;
wire [128*WIDTH-1:0] weight1_3;

wire [32*C_WIDTH-1:0] out_0;
wire [32*C_WIDTH-1:0] out_1;
wire [32*C_WIDTH-1:0] out_2;
wire [32*C_WIDTH-1:0] out_3;
wire [32*C_WIDTH-1:0] out_4;
wire [32*C_WIDTH-1:0] out_5;
wire [32*C_WIDTH-1:0] out_6;
wire [32*C_WIDTH-1:0] out_7;
wire [32*C_WIDTH-1:0] out_8;
wire [32*C_WIDTH-1:0] out_9;
wire [32*C_WIDTH-1:0] out_10;
wire [32*C_WIDTH-1:0] out_11;
wire [32*C_WIDTH-1:0] out_12;
wire [32*C_WIDTH-1:0] out_13;
wire [32*C_WIDTH-1:0] out_14;
wire [32*C_WIDTH-1:0] out_15;
wire [32*C_WIDTH-1:0] out_16;
wire [32*C_WIDTH-1:0] out_17;
wire [32*C_WIDTH-1:0] out_18;
wire [32*C_WIDTH-1:0] out_19;
wire [32*C_WIDTH-1:0] out_20;
wire [32*C_WIDTH-1:0] out_21;
wire [32*C_WIDTH-1:0] out_22;
wire [32*C_WIDTH-1:0] out_23;
wire [32*C_WIDTH-1:0] out_24;
wire [32*C_WIDTH-1:0] out_25;
wire [32*C_WIDTH-1:0] out_26;
wire [32*C_WIDTH-1:0] out_27;
wire [32*C_WIDTH-1:0] out_28;
wire [32*C_WIDTH-1:0] out_29;
wire [32*C_WIDTH-1:0] out_30;
wire [32*C_WIDTH-1:0] out_31;
wire [32*C_WIDTH-1:0] out_32;
wire [32*C_WIDTH-1:0] out_33;
wire [32*C_WIDTH-1:0] out_34;
wire [32*C_WIDTH-1:0] out_35;
wire [32*C_WIDTH-1:0] out_36;
wire [32*C_WIDTH-1:0] out_37;
wire [32*C_WIDTH-1:0] out_38;
wire [32*C_WIDTH-1:0] out_39;
wire [32*C_WIDTH-1:0] out_40;
wire [32*C_WIDTH-1:0] out_41;
wire [32*C_WIDTH-1:0] out_42;
wire [32*C_WIDTH-1:0] out_43;
wire [32*C_WIDTH-1:0] out_44;
wire [32*C_WIDTH-1:0] out_45;
wire [32*C_WIDTH-1:0] out_46;
wire [32*C_WIDTH-1:0] out_47;
wire [32*C_WIDTH-1:0] out_48;
wire [32*C_WIDTH-1:0] out_49;
wire [32*C_WIDTH-1:0] out_50;
wire [32*C_WIDTH-1:0] out_51;
wire [32*C_WIDTH-1:0] out_52;
wire [32*C_WIDTH-1:0] out_53;
wire [32*C_WIDTH-1:0] out_54;
wire [32*C_WIDTH-1:0] out_55;
wire [32*C_WIDTH-1:0] out_56;
wire [32*C_WIDTH-1:0] out_57;
wire [32*C_WIDTH-1:0] out_58;
wire [32*C_WIDTH-1:0] out_59;
wire [32*C_WIDTH-1:0] out_60;
wire [32*C_WIDTH-1:0] out_61;
wire [32*C_WIDTH-1:0] out_62;
wire [32*C_WIDTH-1:0] out_63;
wire [32*C_WIDTH-1:0] out_64;
wire [32*C_WIDTH-1:0] out_65;
wire [32*C_WIDTH-1:0] out_66;
wire [32*C_WIDTH-1:0] out_67;
wire [32*C_WIDTH-1:0] out_68;
wire [32*C_WIDTH-1:0] out_69;
wire [32*C_WIDTH-1:0] out_70;
wire [32*C_WIDTH-1:0] out_71;
wire [32*C_WIDTH-1:0] out_72;
wire [32*C_WIDTH-1:0] out_73;
wire [32*C_WIDTH-1:0] out_74;
wire [32*C_WIDTH-1:0] out_75;
wire [32*C_WIDTH-1:0] out_76;
wire [32*C_WIDTH-1:0] out_77;
wire [32*C_WIDTH-1:0] out_78;
wire [32*C_WIDTH-1:0] out_79;
wire [32*C_WIDTH-1:0] out_80;
wire [32*C_WIDTH-1:0] out_81;
wire [32*C_WIDTH-1:0] out_82;
wire [32*C_WIDTH-1:0] out_83;
wire [32*C_WIDTH-1:0] out_84;
wire [32*C_WIDTH-1:0] out_85;
wire [32*C_WIDTH-1:0] out_86;
wire [32*C_WIDTH-1:0] out_87;
wire [32*C_WIDTH-1:0] out_88;
wire [32*C_WIDTH-1:0] out_89;
wire [32*C_WIDTH-1:0] out_90;
wire [32*C_WIDTH-1:0] out_91;
wire [32*C_WIDTH-1:0] out_92;
wire [32*C_WIDTH-1:0] out_93;
wire [32*C_WIDTH-1:0] out_94;
wire [32*C_WIDTH-1:0] out_95;
wire [32*C_WIDTH-1:0] out_96;
wire [32*C_WIDTH-1:0] out_97;
wire [32*C_WIDTH-1:0] out_98;
wire [32*C_WIDTH-1:0] out_99;
wire [32*C_WIDTH-1:0] out_100;
wire [32*C_WIDTH-1:0] out_101;
wire [32*C_WIDTH-1:0] out_102;
wire [32*C_WIDTH-1:0] out_103;
wire [32*C_WIDTH-1:0] out_104;
wire [32*C_WIDTH-1:0] out_105;
wire [32*C_WIDTH-1:0] out_106;
wire [32*C_WIDTH-1:0] out_107;
wire [32*C_WIDTH-1:0] out_108;
wire [32*C_WIDTH-1:0] out_109;
wire [32*C_WIDTH-1:0] out_110;
wire [32*C_WIDTH-1:0] out_111;
wire [32*C_WIDTH-1:0] out_112;
wire [32*C_WIDTH-1:0] out_113;
wire [32*C_WIDTH-1:0] out_114;
wire [32*C_WIDTH-1:0] out_115;
wire [32*C_WIDTH-1:0] out_116;
wire [32*C_WIDTH-1:0] out_117;
wire [32*C_WIDTH-1:0] out_118;
wire [32*C_WIDTH-1:0] out_119;
wire [32*C_WIDTH-1:0] out_120;
wire [32*C_WIDTH-1:0] out_121;
wire [32*C_WIDTH-1:0] out_122;
wire [32*C_WIDTH-1:0] out_123;
wire [32*C_WIDTH-1:0] out_124;
wire [32*C_WIDTH-1:0] out_125;
wire [32*C_WIDTH-1:0] out_126;
wire [32*C_WIDTH-1:0] out_127;
wire [32*C_WIDTH-1:0] out_128;
wire [32*C_WIDTH-1:0] out_129;
wire [32*C_WIDTH-1:0] out_130;
wire [32*C_WIDTH-1:0] out_131;
wire [32*C_WIDTH-1:0] out_132;
wire [32*C_WIDTH-1:0] out_133;
wire [32*C_WIDTH-1:0] out_134;
wire [32*C_WIDTH-1:0] out_135;
wire [32*C_WIDTH-1:0] out_136;
wire [32*C_WIDTH-1:0] out_137;
wire [32*C_WIDTH-1:0] out_138;
wire [32*C_WIDTH-1:0] out_139;
wire [32*C_WIDTH-1:0] out_140;
wire [32*C_WIDTH-1:0] out_141;
wire [32*C_WIDTH-1:0] out_142;
wire [32*C_WIDTH-1:0] out_143;
wire [32*C_WIDTH-1:0] out_144;
wire [32*C_WIDTH-1:0] out_145;
wire [32*C_WIDTH-1:0] out_146;
wire [32*C_WIDTH-1:0] out_147;
wire [32*C_WIDTH-1:0] out_148;
wire [32*C_WIDTH-1:0] out_149;
wire [32*C_WIDTH-1:0] out_150;
wire [32*C_WIDTH-1:0] out_151;
wire [32*C_WIDTH-1:0] out_152;
wire [32*C_WIDTH-1:0] out_153;
wire [32*C_WIDTH-1:0] out_154;
wire [32*C_WIDTH-1:0] out_155;
wire [32*C_WIDTH-1:0] out_156;
wire [32*C_WIDTH-1:0] out_157;
wire [32*C_WIDTH-1:0] out_158;
wire [32*C_WIDTH-1:0] out_159;
wire [32*C_WIDTH-1:0] out_160;
wire [32*C_WIDTH-1:0] out_161;
wire [32*C_WIDTH-1:0] out_162;
wire [32*C_WIDTH-1:0] out_163;
wire [32*C_WIDTH-1:0] out_164;
wire [32*C_WIDTH-1:0] out_165;
wire [32*C_WIDTH-1:0] out_166;
wire [32*C_WIDTH-1:0] out_167;
wire [32*C_WIDTH-1:0] out_168;
wire [32*C_WIDTH-1:0] out_169;
wire [32*C_WIDTH-1:0] out_170;
wire [32*C_WIDTH-1:0] out_171;
wire [32*C_WIDTH-1:0] out_172;
wire [32*C_WIDTH-1:0] out_173;
wire [32*C_WIDTH-1:0] out_174;
wire [32*C_WIDTH-1:0] out_175;
wire [32*C_WIDTH-1:0] out_176;
wire [32*C_WIDTH-1:0] out_177;
wire [32*C_WIDTH-1:0] out_178;
wire [32*C_WIDTH-1:0] out_179;
wire [32*C_WIDTH-1:0] out_180;
wire [32*C_WIDTH-1:0] out_181;
wire [32*C_WIDTH-1:0] out_182;
wire [32*C_WIDTH-1:0] out_183;
wire [32*C_WIDTH-1:0] out_184;
wire [32*C_WIDTH-1:0] out_185;
wire [32*C_WIDTH-1:0] out_186;
wire [32*C_WIDTH-1:0] out_187;
wire [32*C_WIDTH-1:0] out_188;
wire [32*C_WIDTH-1:0] out_189;
wire [32*C_WIDTH-1:0] out_190;
wire [32*C_WIDTH-1:0] out_191;
wire [32*C_WIDTH-1:0] out_192;
wire [32*C_WIDTH-1:0] out_193;
wire [32*C_WIDTH-1:0] out_194;
wire [32*C_WIDTH-1:0] out_195;
wire [32*C_WIDTH-1:0] out_196;
wire [32*C_WIDTH-1:0] out_197;
wire [32*C_WIDTH-1:0] out_198;
wire [32*C_WIDTH-1:0] out_199;
wire [32*C_WIDTH-1:0] out_200;
wire [32*C_WIDTH-1:0] out_201;
wire [32*C_WIDTH-1:0] out_202;
wire [32*C_WIDTH-1:0] out_203;
wire [32*C_WIDTH-1:0] out_204;
wire [32*C_WIDTH-1:0] out_205;
wire [32*C_WIDTH-1:0] out_206;
wire [32*C_WIDTH-1:0] out_207;
wire [32*C_WIDTH-1:0] out_208;
wire [32*C_WIDTH-1:0] out_209;
wire [32*C_WIDTH-1:0] out_210;
wire [32*C_WIDTH-1:0] out_211;
wire [32*C_WIDTH-1:0] out_212;
wire [32*C_WIDTH-1:0] out_213;
wire [32*C_WIDTH-1:0] out_214;
wire [32*C_WIDTH-1:0] out_215;
wire [32*C_WIDTH-1:0] out_216;
wire [32*C_WIDTH-1:0] out_217;
wire [32*C_WIDTH-1:0] out_218;
wire [32*C_WIDTH-1:0] out_219;
wire [32*C_WIDTH-1:0] out_220;
wire [32*C_WIDTH-1:0] out_221;
wire [32*C_WIDTH-1:0] out_222;
wire [32*C_WIDTH-1:0] out_223;
wire [32*C_WIDTH-1:0] out_224;
wire [32*C_WIDTH-1:0] out_225;
wire [32*C_WIDTH-1:0] out_226;
wire [32*C_WIDTH-1:0] out_227;
wire [32*C_WIDTH-1:0] out_228;
wire [32*C_WIDTH-1:0] out_229;
wire [32*C_WIDTH-1:0] out_230;
wire [32*C_WIDTH-1:0] out_231;
wire [32*C_WIDTH-1:0] out_232;
wire [32*C_WIDTH-1:0] out_233;
wire [32*C_WIDTH-1:0] out_234;
wire [32*C_WIDTH-1:0] out_235;
wire [32*C_WIDTH-1:0] out_236;
wire [32*C_WIDTH-1:0] out_237;
wire [32*C_WIDTH-1:0] out_238;
wire [32*C_WIDTH-1:0] out_239;
wire [32*C_WIDTH-1:0] out_240;
wire [32*C_WIDTH-1:0] out_241;
wire [32*C_WIDTH-1:0] out_242;
wire [32*C_WIDTH-1:0] out_243;
wire [32*C_WIDTH-1:0] out_244;
wire [32*C_WIDTH-1:0] out_245;
wire [32*C_WIDTH-1:0] out_246;
wire [32*C_WIDTH-1:0] out_247;
wire [32*C_WIDTH-1:0] out_248;
wire [32*C_WIDTH-1:0] out_249;
wire [32*C_WIDTH-1:0] out_250;
wire [32*C_WIDTH-1:0] out_251;
wire [32*C_WIDTH-1:0] out_252;
wire [32*C_WIDTH-1:0] out_253;
wire [32*C_WIDTH-1:0] out_254;
wire [32*C_WIDTH-1:0] out_255;
wire [32*C_WIDTH-1:0] out_256;
wire [32*C_WIDTH-1:0] out_257;
wire [32*C_WIDTH-1:0] out_258;
wire [32*C_WIDTH-1:0] out_259;
wire [32*C_WIDTH-1:0] out_260;
wire [32*C_WIDTH-1:0] out_261;
wire [32*C_WIDTH-1:0] out_262;
wire [32*C_WIDTH-1:0] out_263;
wire [32*C_WIDTH-1:0] out_264;
wire [32*C_WIDTH-1:0] out_265;
wire [32*C_WIDTH-1:0] out_266;
wire [32*C_WIDTH-1:0] out_267;
wire [32*C_WIDTH-1:0] out_268;
wire [32*C_WIDTH-1:0] out_269;
wire [32*C_WIDTH-1:0] out_270;
wire [32*C_WIDTH-1:0] out_271;
wire [32*C_WIDTH-1:0] out_272;
wire [32*C_WIDTH-1:0] out_273;
wire [32*C_WIDTH-1:0] out_274;
wire [32*C_WIDTH-1:0] out_275;
wire [32*C_WIDTH-1:0] out_276;
wire [32*C_WIDTH-1:0] out_277;
wire [32*C_WIDTH-1:0] out_278;
wire [32*C_WIDTH-1:0] out_279;
wire [32*C_WIDTH-1:0] out_280;
wire [32*C_WIDTH-1:0] out_281;
wire [32*C_WIDTH-1:0] out_282;
wire [32*C_WIDTH-1:0] out_283;
wire [32*C_WIDTH-1:0] out_284;
wire [32*C_WIDTH-1:0] out_285;
wire [32*C_WIDTH-1:0] out_286;
wire [32*C_WIDTH-1:0] out_287;
wire [32*C_WIDTH-1:0] out_288;
wire [32*C_WIDTH-1:0] out_289;
wire [32*C_WIDTH-1:0] out_290;
wire [32*C_WIDTH-1:0] out_291;
wire [32*C_WIDTH-1:0] out_292;
wire [32*C_WIDTH-1:0] out_293;
wire [32*C_WIDTH-1:0] out_294;
wire [32*C_WIDTH-1:0] out_295;
wire [32*C_WIDTH-1:0] out_296;
wire [32*C_WIDTH-1:0] out_297;
wire [32*C_WIDTH-1:0] out_298;
wire [32*C_WIDTH-1:0] out_299;
wire [32*C_WIDTH-1:0] out_300;
wire [32*C_WIDTH-1:0] out_301;
wire [32*C_WIDTH-1:0] out_302;
wire [32*C_WIDTH-1:0] out_303;
wire [32*C_WIDTH-1:0] out_304;
wire [32*C_WIDTH-1:0] out_305;
wire [32*C_WIDTH-1:0] out_306;
wire [32*C_WIDTH-1:0] out_307;
wire [32*C_WIDTH-1:0] out_308;
wire [32*C_WIDTH-1:0] out_309;
wire [32*C_WIDTH-1:0] out_310;
wire [32*C_WIDTH-1:0] out_311;
wire [32*C_WIDTH-1:0] out_312;
wire [32*C_WIDTH-1:0] out_313;
wire [32*C_WIDTH-1:0] out_314;
wire [32*C_WIDTH-1:0] out_315;
wire [32*C_WIDTH-1:0] out_316;
wire [32*C_WIDTH-1:0] out_317;
wire [32*C_WIDTH-1:0] out_318;
wire [32*C_WIDTH-1:0] out_319;
wire [32*C_WIDTH-1:0] out_320;
wire [32*C_WIDTH-1:0] out_321;
wire [32*C_WIDTH-1:0] out_322;
wire [32*C_WIDTH-1:0] out_323;
wire [32*C_WIDTH-1:0] out_324;
wire [32*C_WIDTH-1:0] out_325;
wire [32*C_WIDTH-1:0] out_326;
wire [32*C_WIDTH-1:0] out_327;
wire [32*C_WIDTH-1:0] out_328;
wire [32*C_WIDTH-1:0] out_329;
wire [32*C_WIDTH-1:0] out_330;
wire [32*C_WIDTH-1:0] out_331;
wire [32*C_WIDTH-1:0] out_332;
wire [32*C_WIDTH-1:0] out_333;
wire [32*C_WIDTH-1:0] out_334;
wire [32*C_WIDTH-1:0] out_335;
wire [32*C_WIDTH-1:0] out_336;
wire [32*C_WIDTH-1:0] out_337;
wire [32*C_WIDTH-1:0] out_338;
wire [32*C_WIDTH-1:0] out_339;
wire [32*C_WIDTH-1:0] out_340;
wire [32*C_WIDTH-1:0] out_341;
wire [32*C_WIDTH-1:0] out_342;
wire [32*C_WIDTH-1:0] out_343;
wire [32*C_WIDTH-1:0] out_344;
wire [32*C_WIDTH-1:0] out_345;
wire [32*C_WIDTH-1:0] out_346;
wire [32*C_WIDTH-1:0] out_347;
wire [32*C_WIDTH-1:0] out_348;
wire [32*C_WIDTH-1:0] out_349;
wire [32*C_WIDTH-1:0] out_350;
wire [32*C_WIDTH-1:0] out_351;
wire [32*C_WIDTH-1:0] out_352;
wire [32*C_WIDTH-1:0] out_353;
wire [32*C_WIDTH-1:0] out_354;
wire [32*C_WIDTH-1:0] out_355;
wire [32*C_WIDTH-1:0] out_356;
wire [32*C_WIDTH-1:0] out_357;
wire [32*C_WIDTH-1:0] out_358;
wire [32*C_WIDTH-1:0] out_359;
wire [32*C_WIDTH-1:0] out_360;
wire [32*C_WIDTH-1:0] out_361;
wire [32*C_WIDTH-1:0] out_362;
wire [32*C_WIDTH-1:0] out_363;
wire [32*C_WIDTH-1:0] out_364;
wire [32*C_WIDTH-1:0] out_365;
wire [32*C_WIDTH-1:0] out_366;
wire [32*C_WIDTH-1:0] out_367;
wire [32*C_WIDTH-1:0] out_368;
wire [32*C_WIDTH-1:0] out_369;
wire [32*C_WIDTH-1:0] out_370;
wire [32*C_WIDTH-1:0] out_371;
wire [32*C_WIDTH-1:0] out_372;
wire [32*C_WIDTH-1:0] out_373;
wire [32*C_WIDTH-1:0] out_374;
wire [32*C_WIDTH-1:0] out_375;
wire [32*C_WIDTH-1:0] out_376;
wire [32*C_WIDTH-1:0] out_377;
wire [32*C_WIDTH-1:0] out_378;
wire [32*C_WIDTH-1:0] out_379;
wire [32*C_WIDTH-1:0] out_380;
wire [32*C_WIDTH-1:0] out_381;
wire [32*C_WIDTH-1:0] out_382;
wire [32*C_WIDTH-1:0] out_383;
wire [32*C_WIDTH-1:0] out_384;
wire [32*C_WIDTH-1:0] out_385;
wire [32*C_WIDTH-1:0] out_386;
wire [32*C_WIDTH-1:0] out_387;
wire [32*C_WIDTH-1:0] out_388;
wire [32*C_WIDTH-1:0] out_389;
wire [32*C_WIDTH-1:0] out_390;
wire [32*C_WIDTH-1:0] out_391;
wire [32*C_WIDTH-1:0] out_392;
wire [32*C_WIDTH-1:0] out_393;
wire [32*C_WIDTH-1:0] out_394;
wire [32*C_WIDTH-1:0] out_395;
wire [32*C_WIDTH-1:0] out_396;
wire [32*C_WIDTH-1:0] out_397;
wire [32*C_WIDTH-1:0] out_398;
wire [32*C_WIDTH-1:0] out_399;
wire [32*C_WIDTH-1:0] out_400;
wire [32*C_WIDTH-1:0] out_401;
wire [32*C_WIDTH-1:0] out_402;
wire [32*C_WIDTH-1:0] out_403;
wire [32*C_WIDTH-1:0] out_404;
wire [32*C_WIDTH-1:0] out_405;
wire [32*C_WIDTH-1:0] out_406;
wire [32*C_WIDTH-1:0] out_407;
wire [32*C_WIDTH-1:0] out_408;
wire [32*C_WIDTH-1:0] out_409;
wire [32*C_WIDTH-1:0] out_410;
wire [32*C_WIDTH-1:0] out_411;
wire [32*C_WIDTH-1:0] out_412;
wire [32*C_WIDTH-1:0] out_413;
wire [32*C_WIDTH-1:0] out_414;
wire [32*C_WIDTH-1:0] out_415;
wire [32*C_WIDTH-1:0] out_416;
wire [32*C_WIDTH-1:0] out_417;
wire [32*C_WIDTH-1:0] out_418;
wire [32*C_WIDTH-1:0] out_419;
wire [32*C_WIDTH-1:0] out_420;
wire [32*C_WIDTH-1:0] out_421;
wire [32*C_WIDTH-1:0] out_422;
wire [32*C_WIDTH-1:0] out_423;
wire [32*C_WIDTH-1:0] out_424;
wire [32*C_WIDTH-1:0] out_425;
wire [32*C_WIDTH-1:0] out_426;
wire [32*C_WIDTH-1:0] out_427;
wire [32*C_WIDTH-1:0] out_428;
wire [32*C_WIDTH-1:0] out_429;
wire [32*C_WIDTH-1:0] out_430;
wire [32*C_WIDTH-1:0] out_431;
wire [32*C_WIDTH-1:0] out_432;
wire [32*C_WIDTH-1:0] out_433;
wire [32*C_WIDTH-1:0] out_434;
wire [32*C_WIDTH-1:0] out_435;
wire [32*C_WIDTH-1:0] out_436;
wire [32*C_WIDTH-1:0] out_437;
wire [32*C_WIDTH-1:0] out_438;
wire [32*C_WIDTH-1:0] out_439;
wire [32*C_WIDTH-1:0] out_440;
wire [32*C_WIDTH-1:0] out_441;
wire [32*C_WIDTH-1:0] out_442;
wire [32*C_WIDTH-1:0] out_443;
wire [32*C_WIDTH-1:0] out_444;
wire [32*C_WIDTH-1:0] out_445;
wire [32*C_WIDTH-1:0] out_446;
wire [32*C_WIDTH-1:0] out_447;
wire [32*C_WIDTH-1:0] out_448;
wire [32*C_WIDTH-1:0] out_449;
wire [32*C_WIDTH-1:0] out_450;
wire [32*C_WIDTH-1:0] out_451;
wire [32*C_WIDTH-1:0] out_452;
wire [32*C_WIDTH-1:0] out_453;
wire [32*C_WIDTH-1:0] out_454;
wire [32*C_WIDTH-1:0] out_455;
wire [32*C_WIDTH-1:0] out_456;
wire [32*C_WIDTH-1:0] out_457;
wire [32*C_WIDTH-1:0] out_458;
wire [32*C_WIDTH-1:0] out_459;
wire [32*C_WIDTH-1:0] out_460;
wire [32*C_WIDTH-1:0] out_461;
wire [32*C_WIDTH-1:0] out_462;
wire [32*C_WIDTH-1:0] out_463;
wire [32*C_WIDTH-1:0] out_464;
wire [32*C_WIDTH-1:0] out_465;
wire [32*C_WIDTH-1:0] out_466;
wire [32*C_WIDTH-1:0] out_467;
wire [32*C_WIDTH-1:0] out_468;
wire [32*C_WIDTH-1:0] out_469;
wire [32*C_WIDTH-1:0] out_470;
wire [32*C_WIDTH-1:0] out_471;
wire [32*C_WIDTH-1:0] out_472;
wire [32*C_WIDTH-1:0] out_473;
wire [32*C_WIDTH-1:0] out_474;
wire [32*C_WIDTH-1:0] out_475;
wire [32*C_WIDTH-1:0] out_476;
wire [32*C_WIDTH-1:0] out_477;
wire [32*C_WIDTH-1:0] out_478;
wire [32*C_WIDTH-1:0] out_479;
wire [32*C_WIDTH-1:0] out_480;
wire [32*C_WIDTH-1:0] out_481;
wire [32*C_WIDTH-1:0] out_482;
wire [32*C_WIDTH-1:0] out_483;
wire [32*C_WIDTH-1:0] out_484;
wire [32*C_WIDTH-1:0] out_485;
wire [32*C_WIDTH-1:0] out_486;
wire [32*C_WIDTH-1:0] out_487;
wire [32*C_WIDTH-1:0] out_488;
wire [32*C_WIDTH-1:0] out_489;
wire [32*C_WIDTH-1:0] out_490;
wire [32*C_WIDTH-1:0] out_491;
wire [32*C_WIDTH-1:0] out_492;
wire [32*C_WIDTH-1:0] out_493;
wire [32*C_WIDTH-1:0] out_494;
wire [32*C_WIDTH-1:0] out_495;
wire [32*C_WIDTH-1:0] out_496;
wire [32*C_WIDTH-1:0] out_497;
wire [32*C_WIDTH-1:0] out_498;
wire [32*C_WIDTH-1:0] out_499;
wire [32*C_WIDTH-1:0] out_500;
wire [32*C_WIDTH-1:0] out_501;
wire [32*C_WIDTH-1:0] out_502;
wire [32*C_WIDTH-1:0] out_503;
wire [32*C_WIDTH-1:0] out_504;
wire [32*C_WIDTH-1:0] out_505;
wire [32*C_WIDTH-1:0] out_506;
wire [32*C_WIDTH-1:0] out_507;
wire [32*C_WIDTH-1:0] out_508;
wire [32*C_WIDTH-1:0] out_509;
wire [32*C_WIDTH-1:0] out_510;
wire [32*C_WIDTH-1:0] out_511;
wire [32*C_WIDTH-1:0] out_512;
wire [32*C_WIDTH-1:0] out_513;
wire [32*C_WIDTH-1:0] out_514;
wire [32*C_WIDTH-1:0] out_515;
wire [32*C_WIDTH-1:0] out_516;
wire [32*C_WIDTH-1:0] out_517;
wire [32*C_WIDTH-1:0] out_518;
wire [32*C_WIDTH-1:0] out_519;
wire [32*C_WIDTH-1:0] out_520;
wire [32*C_WIDTH-1:0] out_521;
wire [32*C_WIDTH-1:0] out_522;
wire [32*C_WIDTH-1:0] out_523;
wire [32*C_WIDTH-1:0] out_524;
wire [32*C_WIDTH-1:0] out_525;
wire [32*C_WIDTH-1:0] out_526;
wire [32*C_WIDTH-1:0] out_527;
wire [32*C_WIDTH-1:0] out_528;
wire [32*C_WIDTH-1:0] out_529;
wire [32*C_WIDTH-1:0] out_530;
wire [32*C_WIDTH-1:0] out_531;
wire [32*C_WIDTH-1:0] out_532;
wire [32*C_WIDTH-1:0] out_533;
wire [32*C_WIDTH-1:0] out_534;
wire [32*C_WIDTH-1:0] out_535;
wire [32*C_WIDTH-1:0] out_536;
wire [32*C_WIDTH-1:0] out_537;
wire [32*C_WIDTH-1:0] out_538;
wire [32*C_WIDTH-1:0] out_539;
wire [32*C_WIDTH-1:0] out_540;
wire [32*C_WIDTH-1:0] out_541;
wire [32*C_WIDTH-1:0] out_542;
wire [32*C_WIDTH-1:0] out_543;
wire [32*C_WIDTH-1:0] out_544;
wire [32*C_WIDTH-1:0] out_545;
wire [32*C_WIDTH-1:0] out_546;
wire [32*C_WIDTH-1:0] out_547;
wire [32*C_WIDTH-1:0] out_548;
wire [32*C_WIDTH-1:0] out_549;
wire [32*C_WIDTH-1:0] out_550;
wire [32*C_WIDTH-1:0] out_551;
wire [32*C_WIDTH-1:0] out_552;
wire [32*C_WIDTH-1:0] out_553;
wire [32*C_WIDTH-1:0] out_554;
wire [32*C_WIDTH-1:0] out_555;
wire [32*C_WIDTH-1:0] out_556;
wire [32*C_WIDTH-1:0] out_557;
wire [32*C_WIDTH-1:0] out_558;
wire [32*C_WIDTH-1:0] out_559;
wire [32*C_WIDTH-1:0] out_560;
wire [32*C_WIDTH-1:0] out_561;
wire [32*C_WIDTH-1:0] out_562;
wire [32*C_WIDTH-1:0] out_563;
wire [32*C_WIDTH-1:0] out_564;
wire [32*C_WIDTH-1:0] out_565;
wire [32*C_WIDTH-1:0] out_566;
wire [32*C_WIDTH-1:0] out_567;
wire [32*C_WIDTH-1:0] out_568;
wire [32*C_WIDTH-1:0] out_569;
wire [32*C_WIDTH-1:0] out_570;
wire [32*C_WIDTH-1:0] out_571;
wire [32*C_WIDTH-1:0] out_572;
wire [32*C_WIDTH-1:0] out_573;
wire [32*C_WIDTH-1:0] out_574;
wire [32*C_WIDTH-1:0] out_575;
wire [32*C_WIDTH-1:0] out_576;
wire [32*C_WIDTH-1:0] out_577;
wire [32*C_WIDTH-1:0] out_578;
wire [32*C_WIDTH-1:0] out_579;
wire [32*C_WIDTH-1:0] out_580;
wire [32*C_WIDTH-1:0] out_581;
wire [32*C_WIDTH-1:0] out_582;
wire [32*C_WIDTH-1:0] out_583;
wire [32*C_WIDTH-1:0] out_584;
wire [32*C_WIDTH-1:0] out_585;
wire [32*C_WIDTH-1:0] out_586;
wire [32*C_WIDTH-1:0] out_587;
wire [32*C_WIDTH-1:0] out_588;
wire [32*C_WIDTH-1:0] out_589;
wire [32*C_WIDTH-1:0] out_590;
wire [32*C_WIDTH-1:0] out_591;
wire [32*C_WIDTH-1:0] out_592;
wire [32*C_WIDTH-1:0] out_593;
wire [32*C_WIDTH-1:0] out_594;
wire [32*C_WIDTH-1:0] out_595;
wire [32*C_WIDTH-1:0] out_596;
wire [32*C_WIDTH-1:0] out_597;
wire [32*C_WIDTH-1:0] out_598;
wire [32*C_WIDTH-1:0] out_599;
wire [32*C_WIDTH-1:0] out_600;
wire [32*C_WIDTH-1:0] out_601;
wire [32*C_WIDTH-1:0] out_602;
wire [32*C_WIDTH-1:0] out_603;
wire [32*C_WIDTH-1:0] out_604;
wire [32*C_WIDTH-1:0] out_605;
wire [32*C_WIDTH-1:0] out_606;
wire [32*C_WIDTH-1:0] out_607;
wire [32*C_WIDTH-1:0] out_608;
wire [32*C_WIDTH-1:0] out_609;
wire [32*C_WIDTH-1:0] out_610;
wire [32*C_WIDTH-1:0] out_611;
wire [32*C_WIDTH-1:0] out_612;
wire [32*C_WIDTH-1:0] out_613;
wire [32*C_WIDTH-1:0] out_614;
wire [32*C_WIDTH-1:0] out_615;
wire [32*C_WIDTH-1:0] out_616;
wire [32*C_WIDTH-1:0] out_617;
wire [32*C_WIDTH-1:0] out_618;
wire [32*C_WIDTH-1:0] out_619;
wire [32*C_WIDTH-1:0] out_620;
wire [32*C_WIDTH-1:0] out_621;
wire [32*C_WIDTH-1:0] out_622;
wire [32*C_WIDTH-1:0] out_623;
wire [32*C_WIDTH-1:0] out_624;
wire [32*C_WIDTH-1:0] out_625;
wire [32*C_WIDTH-1:0] out_626;
wire [32*C_WIDTH-1:0] out_627;
wire [32*C_WIDTH-1:0] out_628;
wire [32*C_WIDTH-1:0] out_629;
wire [32*C_WIDTH-1:0] out_630;
wire [32*C_WIDTH-1:0] out_631;
wire [32*C_WIDTH-1:0] out_632;
wire [32*C_WIDTH-1:0] out_633;
wire [32*C_WIDTH-1:0] out_634;
wire [32*C_WIDTH-1:0] out_635;
wire [32*C_WIDTH-1:0] out_636;
wire [32*C_WIDTH-1:0] out_637;
wire [32*C_WIDTH-1:0] out_638;
wire [32*C_WIDTH-1:0] out_639;
wire [32*C_WIDTH-1:0] out_640;
wire [32*C_WIDTH-1:0] out_641;
wire [32*C_WIDTH-1:0] out_642;
wire [32*C_WIDTH-1:0] out_643;
wire [32*C_WIDTH-1:0] out_644;
wire [32*C_WIDTH-1:0] out_645;
wire [32*C_WIDTH-1:0] out_646;
wire [32*C_WIDTH-1:0] out_647;
wire [32*C_WIDTH-1:0] out_648;
wire [32*C_WIDTH-1:0] out_649;
wire [32*C_WIDTH-1:0] out_650;
wire [32*C_WIDTH-1:0] out_651;
wire [32*C_WIDTH-1:0] out_652;
wire [32*C_WIDTH-1:0] out_653;
wire [32*C_WIDTH-1:0] out_654;
wire [32*C_WIDTH-1:0] out_655;
wire [32*C_WIDTH-1:0] out_656;
wire [32*C_WIDTH-1:0] out_657;
wire [32*C_WIDTH-1:0] out_658;
wire [32*C_WIDTH-1:0] out_659;
wire [32*C_WIDTH-1:0] out_660;
wire [32*C_WIDTH-1:0] out_661;
wire [32*C_WIDTH-1:0] out_662;
wire [32*C_WIDTH-1:0] out_663;
wire [32*C_WIDTH-1:0] out_664;
wire [32*C_WIDTH-1:0] out_665;
wire [32*C_WIDTH-1:0] out_666;
wire [32*C_WIDTH-1:0] out_667;
wire [32*C_WIDTH-1:0] out_668;
wire [32*C_WIDTH-1:0] out_669;
wire [32*C_WIDTH-1:0] out_670;
wire [32*C_WIDTH-1:0] out_671;
wire [32*C_WIDTH-1:0] out_672;
wire [32*C_WIDTH-1:0] out_673;
wire [32*C_WIDTH-1:0] out_674;
wire [32*C_WIDTH-1:0] out_675;
wire [32*C_WIDTH-1:0] out_676;
wire [32*C_WIDTH-1:0] out_677;
wire [32*C_WIDTH-1:0] out_678;
wire [32*C_WIDTH-1:0] out_679;
wire [32*C_WIDTH-1:0] out_680;
wire [32*C_WIDTH-1:0] out_681;
wire [32*C_WIDTH-1:0] out_682;
wire [32*C_WIDTH-1:0] out_683;
wire [32*C_WIDTH-1:0] out_684;
wire [32*C_WIDTH-1:0] out_685;
wire [32*C_WIDTH-1:0] out_686;
wire [32*C_WIDTH-1:0] out_687;
wire [32*C_WIDTH-1:0] out_688;
wire [32*C_WIDTH-1:0] out_689;
wire [32*C_WIDTH-1:0] out_690;
wire [32*C_WIDTH-1:0] out_691;
wire [32*C_WIDTH-1:0] out_692;
wire [32*C_WIDTH-1:0] out_693;
wire [32*C_WIDTH-1:0] out_694;
wire [32*C_WIDTH-1:0] out_695;
wire [32*C_WIDTH-1:0] out_696;
wire [32*C_WIDTH-1:0] out_697;
wire [32*C_WIDTH-1:0] out_698;
wire [32*C_WIDTH-1:0] out_699;
wire [32*C_WIDTH-1:0] out_700;
wire [32*C_WIDTH-1:0] out_701;
wire [32*C_WIDTH-1:0] out_702;
wire [32*C_WIDTH-1:0] out_703;
wire [32*C_WIDTH-1:0] out_704;
wire [32*C_WIDTH-1:0] out_705;
wire [32*C_WIDTH-1:0] out_706;
wire [32*C_WIDTH-1:0] out_707;
wire [32*C_WIDTH-1:0] out_708;
wire [32*C_WIDTH-1:0] out_709;
wire [32*C_WIDTH-1:0] out_710;
wire [32*C_WIDTH-1:0] out_711;
wire [32*C_WIDTH-1:0] out_712;
wire [32*C_WIDTH-1:0] out_713;
wire [32*C_WIDTH-1:0] out_714;
wire [32*C_WIDTH-1:0] out_715;
wire [32*C_WIDTH-1:0] out_716;
wire [32*C_WIDTH-1:0] out_717;
wire [32*C_WIDTH-1:0] out_718;
wire [32*C_WIDTH-1:0] out_719;
wire [32*C_WIDTH-1:0] out_720;
wire [32*C_WIDTH-1:0] out_721;
wire [32*C_WIDTH-1:0] out_722;
wire [32*C_WIDTH-1:0] out_723;
wire [32*C_WIDTH-1:0] out_724;
wire [32*C_WIDTH-1:0] out_725;
wire [32*C_WIDTH-1:0] out_726;
wire [32*C_WIDTH-1:0] out_727;
wire [32*C_WIDTH-1:0] out_728;
wire [32*C_WIDTH-1:0] out_729;
wire [32*C_WIDTH-1:0] out_730;
wire [32*C_WIDTH-1:0] out_731;
wire [32*C_WIDTH-1:0] out_732;
wire [32*C_WIDTH-1:0] out_733;
wire [32*C_WIDTH-1:0] out_734;
wire [32*C_WIDTH-1:0] out_735;
wire [32*C_WIDTH-1:0] out_736;
wire [32*C_WIDTH-1:0] out_737;
wire [32*C_WIDTH-1:0] out_738;
wire [32*C_WIDTH-1:0] out_739;
wire [32*C_WIDTH-1:0] out_740;
wire [32*C_WIDTH-1:0] out_741;
wire [32*C_WIDTH-1:0] out_742;
wire [32*C_WIDTH-1:0] out_743;
wire [32*C_WIDTH-1:0] out_744;
wire [32*C_WIDTH-1:0] out_745;
wire [32*C_WIDTH-1:0] out_746;
wire [32*C_WIDTH-1:0] out_747;
wire [32*C_WIDTH-1:0] out_748;
wire [32*C_WIDTH-1:0] out_749;
wire [32*C_WIDTH-1:0] out_750;
wire [32*C_WIDTH-1:0] out_751;
wire [32*C_WIDTH-1:0] out_752;
wire [32*C_WIDTH-1:0] out_753;
wire [32*C_WIDTH-1:0] out_754;
wire [32*C_WIDTH-1:0] out_755;
wire [32*C_WIDTH-1:0] out_756;
wire [32*C_WIDTH-1:0] out_757;
wire [32*C_WIDTH-1:0] out_758;
wire [32*C_WIDTH-1:0] out_759;
wire [32*C_WIDTH-1:0] out_760;
wire [32*C_WIDTH-1:0] out_761;
wire [32*C_WIDTH-1:0] out_762;
wire [32*C_WIDTH-1:0] out_763;
wire [32*C_WIDTH-1:0] out_764;
wire [32*C_WIDTH-1:0] out_765;
wire [32*C_WIDTH-1:0] out_766;
wire [32*C_WIDTH-1:0] out_767;
wire [32*C_WIDTH-1:0] out_768;
wire [32*C_WIDTH-1:0] out_769;
wire [32*C_WIDTH-1:0] out_770;
wire [32*C_WIDTH-1:0] out_771;
wire [32*C_WIDTH-1:0] out_772;
wire [32*C_WIDTH-1:0] out_773;
wire [32*C_WIDTH-1:0] out_774;
wire [32*C_WIDTH-1:0] out_775;
wire [32*C_WIDTH-1:0] out_776;
wire [32*C_WIDTH-1:0] out_777;
wire [32*C_WIDTH-1:0] out_778;
wire [32*C_WIDTH-1:0] out_779;
wire [32*C_WIDTH-1:0] out_780;
wire [32*C_WIDTH-1:0] out_781;
wire [32*C_WIDTH-1:0] out_782;
wire [32*C_WIDTH-1:0] out_783;
wire [32*C_WIDTH-1:0] out_784;
wire [32*C_WIDTH-1:0] out_785;
wire [32*C_WIDTH-1:0] out_786;
wire [32*C_WIDTH-1:0] out_787;
wire [32*C_WIDTH-1:0] out_788;
wire [32*C_WIDTH-1:0] out_789;
wire [32*C_WIDTH-1:0] out_790;
wire [32*C_WIDTH-1:0] out_791;
wire [32*C_WIDTH-1:0] out_792;
wire [32*C_WIDTH-1:0] out_793;
wire [32*C_WIDTH-1:0] out_794;
wire [32*C_WIDTH-1:0] out_795;
wire [32*C_WIDTH-1:0] out_796;
wire [32*C_WIDTH-1:0] out_797;
wire [32*C_WIDTH-1:0] out_798;
wire [32*C_WIDTH-1:0] out_799;
wire [32*C_WIDTH-1:0] out_800;
wire [32*C_WIDTH-1:0] out_801;
wire [32*C_WIDTH-1:0] out_802;
wire [32*C_WIDTH-1:0] out_803;
wire [32*C_WIDTH-1:0] out_804;
wire [32*C_WIDTH-1:0] out_805;
wire [32*C_WIDTH-1:0] out_806;
wire [32*C_WIDTH-1:0] out_807;
wire [32*C_WIDTH-1:0] out_808;
wire [32*C_WIDTH-1:0] out_809;
wire [32*C_WIDTH-1:0] out_810;
wire [32*C_WIDTH-1:0] out_811;
wire [32*C_WIDTH-1:0] out_812;
wire [32*C_WIDTH-1:0] out_813;
wire [32*C_WIDTH-1:0] out_814;
wire [32*C_WIDTH-1:0] out_815;
wire [32*C_WIDTH-1:0] out_816;
wire [32*C_WIDTH-1:0] out_817;
wire [32*C_WIDTH-1:0] out_818;
wire [32*C_WIDTH-1:0] out_819;
wire [32*C_WIDTH-1:0] out_820;
wire [32*C_WIDTH-1:0] out_821;
wire [32*C_WIDTH-1:0] out_822;
wire [32*C_WIDTH-1:0] out_823;
wire [32*C_WIDTH-1:0] out_824;
wire [32*C_WIDTH-1:0] out_825;
wire [32*C_WIDTH-1:0] out_826;
wire [32*C_WIDTH-1:0] out_827;
wire [32*C_WIDTH-1:0] out_828;
wire [32*C_WIDTH-1:0] out_829;
wire [32*C_WIDTH-1:0] out_830;
wire [32*C_WIDTH-1:0] out_831;
wire [32*C_WIDTH-1:0] out_832;
wire [32*C_WIDTH-1:0] out_833;
wire [32*C_WIDTH-1:0] out_834;
wire [32*C_WIDTH-1:0] out_835;
wire [32*C_WIDTH-1:0] out_836;
wire [32*C_WIDTH-1:0] out_837;
wire [32*C_WIDTH-1:0] out_838;
wire [32*C_WIDTH-1:0] out_839;
wire [32*C_WIDTH-1:0] out_840;
wire [32*C_WIDTH-1:0] out_841;
wire [32*C_WIDTH-1:0] out_842;
wire [32*C_WIDTH-1:0] out_843;
wire [32*C_WIDTH-1:0] out_844;
wire [32*C_WIDTH-1:0] out_845;
wire [32*C_WIDTH-1:0] out_846;
wire [32*C_WIDTH-1:0] out_847;
wire [32*C_WIDTH-1:0] out_848;
wire [32*C_WIDTH-1:0] out_849;
wire [32*C_WIDTH-1:0] out_850;
wire [32*C_WIDTH-1:0] out_851;
wire [32*C_WIDTH-1:0] out_852;
wire [32*C_WIDTH-1:0] out_853;
wire [32*C_WIDTH-1:0] out_854;
wire [32*C_WIDTH-1:0] out_855;
wire [32*C_WIDTH-1:0] out_856;
wire [32*C_WIDTH-1:0] out_857;
wire [32*C_WIDTH-1:0] out_858;
wire [32*C_WIDTH-1:0] out_859;
wire [32*C_WIDTH-1:0] out_860;
wire [32*C_WIDTH-1:0] out_861;
wire [32*C_WIDTH-1:0] out_862;
wire [32*C_WIDTH-1:0] out_863;
wire [32*C_WIDTH-1:0] out_864;
wire [32*C_WIDTH-1:0] out_865;
wire [32*C_WIDTH-1:0] out_866;
wire [32*C_WIDTH-1:0] out_867;
wire [32*C_WIDTH-1:0] out_868;
wire [32*C_WIDTH-1:0] out_869;
wire [32*C_WIDTH-1:0] out_870;
wire [32*C_WIDTH-1:0] out_871;
wire [32*C_WIDTH-1:0] out_872;
wire [32*C_WIDTH-1:0] out_873;
wire [32*C_WIDTH-1:0] out_874;
wire [32*C_WIDTH-1:0] out_875;
wire [32*C_WIDTH-1:0] out_876;
wire [32*C_WIDTH-1:0] out_877;
wire [32*C_WIDTH-1:0] out_878;
wire [32*C_WIDTH-1:0] out_879;
wire [32*C_WIDTH-1:0] out_880;
wire [32*C_WIDTH-1:0] out_881;
wire [32*C_WIDTH-1:0] out_882;
wire [32*C_WIDTH-1:0] out_883;
wire [32*C_WIDTH-1:0] out_884;
wire [32*C_WIDTH-1:0] out_885;
wire [32*C_WIDTH-1:0] out_886;
wire [32*C_WIDTH-1:0] out_887;
wire [32*C_WIDTH-1:0] out_888;
wire [32*C_WIDTH-1:0] out_889;
wire [32*C_WIDTH-1:0] out_890;
wire [32*C_WIDTH-1:0] out_891;
wire [32*C_WIDTH-1:0] out_892;
wire [32*C_WIDTH-1:0] out_893;
wire [32*C_WIDTH-1:0] out_894;
wire [32*C_WIDTH-1:0] out_895;
wire [32*C_WIDTH-1:0] out_896;
wire [32*C_WIDTH-1:0] out_897;
wire [32*C_WIDTH-1:0] out_898;
wire [32*C_WIDTH-1:0] out_899;
wire [32*C_WIDTH-1:0] out_900;
wire [32*C_WIDTH-1:0] out_901;
wire [32*C_WIDTH-1:0] out_902;
wire [32*C_WIDTH-1:0] out_903;
wire [32*C_WIDTH-1:0] out_904;
wire [32*C_WIDTH-1:0] out_905;
wire [32*C_WIDTH-1:0] out_906;
wire [32*C_WIDTH-1:0] out_907;
wire [32*C_WIDTH-1:0] out_908;
wire [32*C_WIDTH-1:0] out_909;
wire [32*C_WIDTH-1:0] out_910;
wire [32*C_WIDTH-1:0] out_911;
wire [32*C_WIDTH-1:0] out_912;
wire [32*C_WIDTH-1:0] out_913;
wire [32*C_WIDTH-1:0] out_914;
wire [32*C_WIDTH-1:0] out_915;
wire [32*C_WIDTH-1:0] out_916;
wire [32*C_WIDTH-1:0] out_917;
wire [32*C_WIDTH-1:0] out_918;
wire [32*C_WIDTH-1:0] out_919;
wire [32*C_WIDTH-1:0] out_920;
wire [32*C_WIDTH-1:0] out_921;
wire [32*C_WIDTH-1:0] out_922;
wire [32*C_WIDTH-1:0] out_923;
wire [32*C_WIDTH-1:0] out_924;
wire [32*C_WIDTH-1:0] out_925;
wire [32*C_WIDTH-1:0] out_926;
wire [32*C_WIDTH-1:0] out_927;
wire [32*C_WIDTH-1:0] out_928;
wire [32*C_WIDTH-1:0] out_929;
wire [32*C_WIDTH-1:0] out_930;
wire [32*C_WIDTH-1:0] out_931;
wire [32*C_WIDTH-1:0] out_932;
wire [32*C_WIDTH-1:0] out_933;
wire [32*C_WIDTH-1:0] out_934;
wire [32*C_WIDTH-1:0] out_935;
wire [32*C_WIDTH-1:0] out_936;
wire [32*C_WIDTH-1:0] out_937;
wire [32*C_WIDTH-1:0] out_938;
wire [32*C_WIDTH-1:0] out_939;
wire [32*C_WIDTH-1:0] out_940;
wire [32*C_WIDTH-1:0] out_941;
wire [32*C_WIDTH-1:0] out_942;
wire [32*C_WIDTH-1:0] out_943;
wire [32*C_WIDTH-1:0] out_944;
wire [32*C_WIDTH-1:0] out_945;
wire [32*C_WIDTH-1:0] out_946;
wire [32*C_WIDTH-1:0] out_947;
wire [32*C_WIDTH-1:0] out_948;
wire [32*C_WIDTH-1:0] out_949;
wire [32*C_WIDTH-1:0] out_950;
wire [32*C_WIDTH-1:0] out_951;
wire [32*C_WIDTH-1:0] out_952;
wire [32*C_WIDTH-1:0] out_953;
wire [32*C_WIDTH-1:0] out_954;
wire [32*C_WIDTH-1:0] out_955;
wire [32*C_WIDTH-1:0] out_956;
wire [32*C_WIDTH-1:0] out_957;
wire [32*C_WIDTH-1:0] out_958;
wire [32*C_WIDTH-1:0] out_959;
wire [32*C_WIDTH-1:0] out_960;
wire [32*C_WIDTH-1:0] out_961;
wire [32*C_WIDTH-1:0] out_962;
wire [32*C_WIDTH-1:0] out_963;
wire [32*C_WIDTH-1:0] out_964;
wire [32*C_WIDTH-1:0] out_965;
wire [32*C_WIDTH-1:0] out_966;
wire [32*C_WIDTH-1:0] out_967;
wire [32*C_WIDTH-1:0] out_968;
wire [32*C_WIDTH-1:0] out_969;
wire [32*C_WIDTH-1:0] out_970;
wire [32*C_WIDTH-1:0] out_971;
wire [32*C_WIDTH-1:0] out_972;
wire [32*C_WIDTH-1:0] out_973;
wire [32*C_WIDTH-1:0] out_974;
wire [32*C_WIDTH-1:0] out_975;
wire [32*C_WIDTH-1:0] out_976;
wire [32*C_WIDTH-1:0] out_977;
wire [32*C_WIDTH-1:0] out_978;
wire [32*C_WIDTH-1:0] out_979;
wire [32*C_WIDTH-1:0] out_980;
wire [32*C_WIDTH-1:0] out_981;
wire [32*C_WIDTH-1:0] out_982;
wire [32*C_WIDTH-1:0] out_983;
wire [32*C_WIDTH-1:0] out_984;
wire [32*C_WIDTH-1:0] out_985;
wire [32*C_WIDTH-1:0] out_986;
wire [32*C_WIDTH-1:0] out_987;
wire [32*C_WIDTH-1:0] out_988;
wire [32*C_WIDTH-1:0] out_989;
wire [32*C_WIDTH-1:0] out_990;
wire [32*C_WIDTH-1:0] out_991;
wire [32*C_WIDTH-1:0] out_992;
wire [32*C_WIDTH-1:0] out_993;
wire [32*C_WIDTH-1:0] out_994;
wire [32*C_WIDTH-1:0] out_995;
wire [32*C_WIDTH-1:0] out_996;
wire [32*C_WIDTH-1:0] out_997;
wire [32*C_WIDTH-1:0] out_998;
wire [32*C_WIDTH-1:0] out_999;
wire [32*C_WIDTH-1:0] out_1000;
wire [32*C_WIDTH-1:0] out_1001;
wire [32*C_WIDTH-1:0] out_1002;
wire [32*C_WIDTH-1:0] out_1003;
wire [32*C_WIDTH-1:0] out_1004;
wire [32*C_WIDTH-1:0] out_1005;
wire [32*C_WIDTH-1:0] out_1006;
wire [32*C_WIDTH-1:0] out_1007;
wire [32*C_WIDTH-1:0] out_1008;
wire [32*C_WIDTH-1:0] out_1009;
wire [32*C_WIDTH-1:0] out_1010;
wire [32*C_WIDTH-1:0] out_1011;
wire [32*C_WIDTH-1:0] out_1012;
wire [32*C_WIDTH-1:0] out_1013;
wire [32*C_WIDTH-1:0] out_1014;
wire [32*C_WIDTH-1:0] out_1015;
wire [32*C_WIDTH-1:0] out_1016;
wire [32*C_WIDTH-1:0] out_1017;
wire [32*C_WIDTH-1:0] out_1018;
wire [32*C_WIDTH-1:0] out_1019;
wire [32*C_WIDTH-1:0] out_1020;
wire [32*C_WIDTH-1:0] out_1021;
wire [32*C_WIDTH-1:0] out_1022;
wire [32*C_WIDTH-1:0] out_1023;
wire [32*C_WIDTH-1:0] out_1024;
wire [32*C_WIDTH-1:0] out_1025;
wire [32*C_WIDTH-1:0] out_1026;
wire [32*C_WIDTH-1:0] out_1027;
wire [32*C_WIDTH-1:0] out_1028;
wire [32*C_WIDTH-1:0] out_1029;
wire [32*C_WIDTH-1:0] out_1030;
wire [32*C_WIDTH-1:0] out_1031;
wire [32*C_WIDTH-1:0] out_1032;
wire [32*C_WIDTH-1:0] out_1033;
wire [32*C_WIDTH-1:0] out_1034;
wire [32*C_WIDTH-1:0] out_1035;
wire [32*C_WIDTH-1:0] out_1036;
wire [32*C_WIDTH-1:0] out_1037;
wire [32*C_WIDTH-1:0] out_1038;
wire [32*C_WIDTH-1:0] out_1039;
wire [32*C_WIDTH-1:0] out_1040;
wire [32*C_WIDTH-1:0] out_1041;
wire [32*C_WIDTH-1:0] out_1042;
wire [32*C_WIDTH-1:0] out_1043;
wire [32*C_WIDTH-1:0] out_1044;
wire [32*C_WIDTH-1:0] out_1045;
wire [32*C_WIDTH-1:0] out_1046;
wire [32*C_WIDTH-1:0] out_1047;
wire [32*C_WIDTH-1:0] out_1048;
wire [32*C_WIDTH-1:0] out_1049;
wire [32*C_WIDTH-1:0] out_1050;
wire [32*C_WIDTH-1:0] out_1051;
wire [32*C_WIDTH-1:0] out_1052;
wire [32*C_WIDTH-1:0] out_1053;
wire [32*C_WIDTH-1:0] out_1054;
wire [32*C_WIDTH-1:0] out_1055;
wire [32*C_WIDTH-1:0] out_1056;
wire [32*C_WIDTH-1:0] out_1057;
wire [32*C_WIDTH-1:0] out_1058;
wire [32*C_WIDTH-1:0] out_1059;
wire [32*C_WIDTH-1:0] out_1060;
wire [32*C_WIDTH-1:0] out_1061;
wire [32*C_WIDTH-1:0] out_1062;
wire [32*C_WIDTH-1:0] out_1063;
wire [32*C_WIDTH-1:0] out_1064;
wire [32*C_WIDTH-1:0] out_1065;
wire [32*C_WIDTH-1:0] out_1066;
wire [32*C_WIDTH-1:0] out_1067;
wire [32*C_WIDTH-1:0] out_1068;
wire [32*C_WIDTH-1:0] out_1069;
wire [32*C_WIDTH-1:0] out_1070;
wire [32*C_WIDTH-1:0] out_1071;
wire [32*C_WIDTH-1:0] out_1072;
wire [32*C_WIDTH-1:0] out_1073;
wire [32*C_WIDTH-1:0] out_1074;
wire [32*C_WIDTH-1:0] out_1075;
wire [32*C_WIDTH-1:0] out_1076;
wire [32*C_WIDTH-1:0] out_1077;
wire [32*C_WIDTH-1:0] out_1078;
wire [32*C_WIDTH-1:0] out_1079;
wire [32*C_WIDTH-1:0] out_1080;
wire [32*C_WIDTH-1:0] out_1081;
wire [32*C_WIDTH-1:0] out_1082;
wire [32*C_WIDTH-1:0] out_1083;
wire [32*C_WIDTH-1:0] out_1084;
wire [32*C_WIDTH-1:0] out_1085;
wire [32*C_WIDTH-1:0] out_1086;
wire [32*C_WIDTH-1:0] out_1087;
wire [32*C_WIDTH-1:0] out_1088;
wire [32*C_WIDTH-1:0] out_1089;
wire [32*C_WIDTH-1:0] out_1090;
wire [32*C_WIDTH-1:0] out_1091;
wire [32*C_WIDTH-1:0] out_1092;
wire [32*C_WIDTH-1:0] out_1093;
wire [32*C_WIDTH-1:0] out_1094;
wire [32*C_WIDTH-1:0] out_1095;
wire [32*C_WIDTH-1:0] out_1096;
wire [32*C_WIDTH-1:0] out_1097;
wire [32*C_WIDTH-1:0] out_1098;
wire [32*C_WIDTH-1:0] out_1099;
wire [32*C_WIDTH-1:0] out_1100;
wire [32*C_WIDTH-1:0] out_1101;
wire [32*C_WIDTH-1:0] out_1102;
wire [32*C_WIDTH-1:0] out_1103;
wire [32*C_WIDTH-1:0] out_1104;
wire [32*C_WIDTH-1:0] out_1105;
wire [32*C_WIDTH-1:0] out_1106;
wire [32*C_WIDTH-1:0] out_1107;
wire [32*C_WIDTH-1:0] out_1108;
wire [32*C_WIDTH-1:0] out_1109;
wire [32*C_WIDTH-1:0] out_1110;
wire [32*C_WIDTH-1:0] out_1111;
wire [32*C_WIDTH-1:0] out_1112;
wire [32*C_WIDTH-1:0] out_1113;
wire [32*C_WIDTH-1:0] out_1114;
wire [32*C_WIDTH-1:0] out_1115;
wire [32*C_WIDTH-1:0] out_1116;
wire [32*C_WIDTH-1:0] out_1117;
wire [32*C_WIDTH-1:0] out_1118;
wire [32*C_WIDTH-1:0] out_1119;
wire [32*C_WIDTH-1:0] out_1120;
wire [32*C_WIDTH-1:0] out_1121;
wire [32*C_WIDTH-1:0] out_1122;
wire [32*C_WIDTH-1:0] out_1123;
wire [32*C_WIDTH-1:0] out_1124;
wire [32*C_WIDTH-1:0] out_1125;
wire [32*C_WIDTH-1:0] out_1126;
wire [32*C_WIDTH-1:0] out_1127;
wire [32*C_WIDTH-1:0] out_1128;
wire [32*C_WIDTH-1:0] out_1129;
wire [32*C_WIDTH-1:0] out_1130;
wire [32*C_WIDTH-1:0] out_1131;
wire [32*C_WIDTH-1:0] out_1132;
wire [32*C_WIDTH-1:0] out_1133;
wire [32*C_WIDTH-1:0] out_1134;
wire [32*C_WIDTH-1:0] out_1135;
wire [32*C_WIDTH-1:0] out_1136;
wire [32*C_WIDTH-1:0] out_1137;
wire [32*C_WIDTH-1:0] out_1138;
wire [32*C_WIDTH-1:0] out_1139;
wire [32*C_WIDTH-1:0] out_1140;
wire [32*C_WIDTH-1:0] out_1141;
wire [32*C_WIDTH-1:0] out_1142;
wire [32*C_WIDTH-1:0] out_1143;
wire [32*C_WIDTH-1:0] out_1144;
wire [32*C_WIDTH-1:0] out_1145;
wire [32*C_WIDTH-1:0] out_1146;
wire [32*C_WIDTH-1:0] out_1147;
wire [32*C_WIDTH-1:0] out_1148;
wire [32*C_WIDTH-1:0] out_1149;
wire [32*C_WIDTH-1:0] out_1150;
wire [32*C_WIDTH-1:0] out_1151;
wire [32*C_WIDTH-1:0] out_1152;
wire [32*C_WIDTH-1:0] out_1153;
wire [32*C_WIDTH-1:0] out_1154;
wire [32*C_WIDTH-1:0] out_1155;
wire [32*C_WIDTH-1:0] out_1156;
wire [32*C_WIDTH-1:0] out_1157;
wire [32*C_WIDTH-1:0] out_1158;
wire [32*C_WIDTH-1:0] out_1159;
wire [32*C_WIDTH-1:0] out_1160;
wire [32*C_WIDTH-1:0] out_1161;
wire [32*C_WIDTH-1:0] out_1162;
wire [32*C_WIDTH-1:0] out_1163;
wire [32*C_WIDTH-1:0] out_1164;
wire [32*C_WIDTH-1:0] out_1165;
wire [32*C_WIDTH-1:0] out_1166;
wire [32*C_WIDTH-1:0] out_1167;
wire [32*C_WIDTH-1:0] out_1168;
wire [32*C_WIDTH-1:0] out_1169;
wire [32*C_WIDTH-1:0] out_1170;
wire [32*C_WIDTH-1:0] out_1171;
wire [32*C_WIDTH-1:0] out_1172;
wire [32*C_WIDTH-1:0] out_1173;
wire [32*C_WIDTH-1:0] out_1174;
wire [32*C_WIDTH-1:0] out_1175;
wire [32*C_WIDTH-1:0] out_1176;
wire [32*C_WIDTH-1:0] out_1177;
wire [32*C_WIDTH-1:0] out_1178;
wire [32*C_WIDTH-1:0] out_1179;
wire [32*C_WIDTH-1:0] out_1180;
wire [32*C_WIDTH-1:0] out_1181;
wire [32*C_WIDTH-1:0] out_1182;
wire [32*C_WIDTH-1:0] out_1183;
wire [32*C_WIDTH-1:0] out_1184;
wire [32*C_WIDTH-1:0] out_1185;
wire [32*C_WIDTH-1:0] out_1186;
wire [32*C_WIDTH-1:0] out_1187;
wire [32*C_WIDTH-1:0] out_1188;
wire [32*C_WIDTH-1:0] out_1189;
wire [32*C_WIDTH-1:0] out_1190;
wire [32*C_WIDTH-1:0] out_1191;
wire [32*C_WIDTH-1:0] out_1192;
wire [32*C_WIDTH-1:0] out_1193;
wire [32*C_WIDTH-1:0] out_1194;
wire [32*C_WIDTH-1:0] out_1195;
wire [32*C_WIDTH-1:0] out_1196;
wire [32*C_WIDTH-1:0] out_1197;
wire [32*C_WIDTH-1:0] out_1198;
wire [32*C_WIDTH-1:0] out_1199;
wire [32*C_WIDTH-1:0] out_1200;
wire [32*C_WIDTH-1:0] out_1201;
wire [32*C_WIDTH-1:0] out_1202;
wire [32*C_WIDTH-1:0] out_1203;
wire [32*C_WIDTH-1:0] out_1204;
wire [32*C_WIDTH-1:0] out_1205;
wire [32*C_WIDTH-1:0] out_1206;
wire [32*C_WIDTH-1:0] out_1207;
wire [32*C_WIDTH-1:0] out_1208;
wire [32*C_WIDTH-1:0] out_1209;
wire [32*C_WIDTH-1:0] out_1210;
wire [32*C_WIDTH-1:0] out_1211;
wire [32*C_WIDTH-1:0] out_1212;
wire [32*C_WIDTH-1:0] out_1213;
wire [32*C_WIDTH-1:0] out_1214;
wire [32*C_WIDTH-1:0] out_1215;
wire [32*C_WIDTH-1:0] out_1216;
wire [32*C_WIDTH-1:0] out_1217;
wire [32*C_WIDTH-1:0] out_1218;
wire [32*C_WIDTH-1:0] out_1219;
wire [32*C_WIDTH-1:0] out_1220;
wire [32*C_WIDTH-1:0] out_1221;
wire [32*C_WIDTH-1:0] out_1222;
wire [32*C_WIDTH-1:0] out_1223;
wire [32*C_WIDTH-1:0] out_1224;
wire [32*C_WIDTH-1:0] out_1225;
wire [32*C_WIDTH-1:0] out_1226;
wire [32*C_WIDTH-1:0] out_1227;
wire [32*C_WIDTH-1:0] out_1228;
wire [32*C_WIDTH-1:0] out_1229;
wire [32*C_WIDTH-1:0] out_1230;
wire [32*C_WIDTH-1:0] out_1231;
wire [32*C_WIDTH-1:0] out_1232;
wire [32*C_WIDTH-1:0] out_1233;
wire [32*C_WIDTH-1:0] out_1234;
wire [32*C_WIDTH-1:0] out_1235;
wire [32*C_WIDTH-1:0] out_1236;
wire [32*C_WIDTH-1:0] out_1237;
wire [32*C_WIDTH-1:0] out_1238;
wire [32*C_WIDTH-1:0] out_1239;
wire [32*C_WIDTH-1:0] out_1240;
wire [32*C_WIDTH-1:0] out_1241;
wire [32*C_WIDTH-1:0] out_1242;
wire [32*C_WIDTH-1:0] out_1243;
wire [32*C_WIDTH-1:0] out_1244;
wire [32*C_WIDTH-1:0] out_1245;
wire [32*C_WIDTH-1:0] out_1246;
wire [32*C_WIDTH-1:0] out_1247;
wire [32*C_WIDTH-1:0] out_1248;
wire [32*C_WIDTH-1:0] out_1249;
wire [32*C_WIDTH-1:0] out_1250;
wire [32*C_WIDTH-1:0] out_1251;
wire [32*C_WIDTH-1:0] out_1252;
wire [32*C_WIDTH-1:0] out_1253;
wire [32*C_WIDTH-1:0] out_1254;
wire [32*C_WIDTH-1:0] out_1255;
wire [32*C_WIDTH-1:0] out_1256;
wire [32*C_WIDTH-1:0] out_1257;
wire [32*C_WIDTH-1:0] out_1258;
wire [32*C_WIDTH-1:0] out_1259;
wire [32*C_WIDTH-1:0] out_1260;
wire [32*C_WIDTH-1:0] out_1261;
wire [32*C_WIDTH-1:0] out_1262;
wire [32*C_WIDTH-1:0] out_1263;
wire [32*C_WIDTH-1:0] out_1264;
wire [32*C_WIDTH-1:0] out_1265;
wire [32*C_WIDTH-1:0] out_1266;
wire [32*C_WIDTH-1:0] out_1267;
wire [32*C_WIDTH-1:0] out_1268;
wire [32*C_WIDTH-1:0] out_1269;
wire [32*C_WIDTH-1:0] out_1270;
wire [32*C_WIDTH-1:0] out_1271;
wire [32*C_WIDTH-1:0] out_1272;
wire [32*C_WIDTH-1:0] out_1273;
wire [32*C_WIDTH-1:0] out_1274;
wire [32*C_WIDTH-1:0] out_1275;
wire [32*C_WIDTH-1:0] out_1276;
wire [32*C_WIDTH-1:0] out_1277;
wire [32*C_WIDTH-1:0] out_1278;
wire [32*C_WIDTH-1:0] out_1279;
wire [32*C_WIDTH-1:0] out_1280;
wire [32*C_WIDTH-1:0] out_1281;
wire [32*C_WIDTH-1:0] out_1282;
wire [32*C_WIDTH-1:0] out_1283;
wire [32*C_WIDTH-1:0] out_1284;
wire [32*C_WIDTH-1:0] out_1285;
wire [32*C_WIDTH-1:0] out_1286;
wire [32*C_WIDTH-1:0] out_1287;
wire [32*C_WIDTH-1:0] out_1288;
wire [32*C_WIDTH-1:0] out_1289;
wire [32*C_WIDTH-1:0] out_1290;
wire [32*C_WIDTH-1:0] out_1291;
wire [32*C_WIDTH-1:0] out_1292;
wire [32*C_WIDTH-1:0] out_1293;
wire [32*C_WIDTH-1:0] out_1294;
wire [32*C_WIDTH-1:0] out_1295;
wire [32*C_WIDTH-1:0] out_1296;
wire [32*C_WIDTH-1:0] out_1297;
wire [32*C_WIDTH-1:0] out_1298;
wire [32*C_WIDTH-1:0] out_1299;
wire [32*C_WIDTH-1:0] out_1300;
wire [32*C_WIDTH-1:0] out_1301;
wire [32*C_WIDTH-1:0] out_1302;
wire [32*C_WIDTH-1:0] out_1303;
wire [32*C_WIDTH-1:0] out_1304;
wire [32*C_WIDTH-1:0] out_1305;
wire [32*C_WIDTH-1:0] out_1306;
wire [32*C_WIDTH-1:0] out_1307;
wire [32*C_WIDTH-1:0] out_1308;
wire [32*C_WIDTH-1:0] out_1309;
wire [32*C_WIDTH-1:0] out_1310;
wire [32*C_WIDTH-1:0] out_1311;
wire [32*C_WIDTH-1:0] out_1312;
wire [32*C_WIDTH-1:0] out_1313;
wire [32*C_WIDTH-1:0] out_1314;
wire [32*C_WIDTH-1:0] out_1315;
wire [32*C_WIDTH-1:0] out_1316;
wire [32*C_WIDTH-1:0] out_1317;
wire [32*C_WIDTH-1:0] out_1318;
wire [32*C_WIDTH-1:0] out_1319;
wire [32*C_WIDTH-1:0] out_1320;
wire [32*C_WIDTH-1:0] out_1321;
wire [32*C_WIDTH-1:0] out_1322;
wire [32*C_WIDTH-1:0] out_1323;
wire [32*C_WIDTH-1:0] out_1324;
wire [32*C_WIDTH-1:0] out_1325;
wire [32*C_WIDTH-1:0] out_1326;
wire [32*C_WIDTH-1:0] out_1327;
wire [32*C_WIDTH-1:0] out_1328;
wire [32*C_WIDTH-1:0] out_1329;
wire [32*C_WIDTH-1:0] out_1330;
wire [32*C_WIDTH-1:0] out_1331;
wire [32*C_WIDTH-1:0] out_1332;
wire [32*C_WIDTH-1:0] out_1333;
wire [32*C_WIDTH-1:0] out_1334;
wire [32*C_WIDTH-1:0] out_1335;
wire [32*C_WIDTH-1:0] out_1336;
wire [32*C_WIDTH-1:0] out_1337;
wire [32*C_WIDTH-1:0] out_1338;
wire [32*C_WIDTH-1:0] out_1339;
wire [32*C_WIDTH-1:0] out_1340;
wire [32*C_WIDTH-1:0] out_1341;
wire [32*C_WIDTH-1:0] out_1342;
wire [32*C_WIDTH-1:0] out_1343;
wire [32*C_WIDTH-1:0] out_1344;
wire [32*C_WIDTH-1:0] out_1345;
wire [32*C_WIDTH-1:0] out_1346;
wire [32*C_WIDTH-1:0] out_1347;
wire [32*C_WIDTH-1:0] out_1348;
wire [32*C_WIDTH-1:0] out_1349;
wire [32*C_WIDTH-1:0] out_1350;
wire [32*C_WIDTH-1:0] out_1351;
wire [32*C_WIDTH-1:0] out_1352;
wire [32*C_WIDTH-1:0] out_1353;
wire [32*C_WIDTH-1:0] out_1354;
wire [32*C_WIDTH-1:0] out_1355;
wire [32*C_WIDTH-1:0] out_1356;
wire [32*C_WIDTH-1:0] out_1357;
wire [32*C_WIDTH-1:0] out_1358;
wire [32*C_WIDTH-1:0] out_1359;
wire [32*C_WIDTH-1:0] out_1360;
wire [32*C_WIDTH-1:0] out_1361;
wire [32*C_WIDTH-1:0] out_1362;
wire [32*C_WIDTH-1:0] out_1363;
wire [32*C_WIDTH-1:0] out_1364;
wire [32*C_WIDTH-1:0] out_1365;
wire [32*C_WIDTH-1:0] out_1366;
wire [32*C_WIDTH-1:0] out_1367;
wire [32*C_WIDTH-1:0] out_1368;
wire [32*C_WIDTH-1:0] out_1369;
wire [32*C_WIDTH-1:0] out_1370;
wire [32*C_WIDTH-1:0] out_1371;
wire [32*C_WIDTH-1:0] out_1372;
wire [32*C_WIDTH-1:0] out_1373;
wire [32*C_WIDTH-1:0] out_1374;
wire [32*C_WIDTH-1:0] out_1375;
wire [32*C_WIDTH-1:0] out_1376;
wire [32*C_WIDTH-1:0] out_1377;
wire [32*C_WIDTH-1:0] out_1378;
wire [32*C_WIDTH-1:0] out_1379;
wire [32*C_WIDTH-1:0] out_1380;
wire [32*C_WIDTH-1:0] out_1381;
wire [32*C_WIDTH-1:0] out_1382;
wire [32*C_WIDTH-1:0] out_1383;
wire [32*C_WIDTH-1:0] out_1384;
wire [32*C_WIDTH-1:0] out_1385;
wire [32*C_WIDTH-1:0] out_1386;
wire [32*C_WIDTH-1:0] out_1387;
wire [32*C_WIDTH-1:0] out_1388;
wire [32*C_WIDTH-1:0] out_1389;
wire [32*C_WIDTH-1:0] out_1390;
wire [32*C_WIDTH-1:0] out_1391;
wire [32*C_WIDTH-1:0] out_1392;
wire [32*C_WIDTH-1:0] out_1393;
wire [32*C_WIDTH-1:0] out_1394;
wire [32*C_WIDTH-1:0] out_1395;
wire [32*C_WIDTH-1:0] out_1396;
wire [32*C_WIDTH-1:0] out_1397;
wire [32*C_WIDTH-1:0] out_1398;
wire [32*C_WIDTH-1:0] out_1399;
wire [32*C_WIDTH-1:0] out_1400;
wire [32*C_WIDTH-1:0] out_1401;
wire [32*C_WIDTH-1:0] out_1402;
wire [32*C_WIDTH-1:0] out_1403;
wire [32*C_WIDTH-1:0] out_1404;
wire [32*C_WIDTH-1:0] out_1405;
wire [32*C_WIDTH-1:0] out_1406;
wire [32*C_WIDTH-1:0] out_1407;
wire [32*C_WIDTH-1:0] out_1408;
wire [32*C_WIDTH-1:0] out_1409;
wire [32*C_WIDTH-1:0] out_1410;
wire [32*C_WIDTH-1:0] out_1411;
wire [32*C_WIDTH-1:0] out_1412;
wire [32*C_WIDTH-1:0] out_1413;
wire [32*C_WIDTH-1:0] out_1414;
wire [32*C_WIDTH-1:0] out_1415;
wire [32*C_WIDTH-1:0] out_1416;
wire [32*C_WIDTH-1:0] out_1417;
wire [32*C_WIDTH-1:0] out_1418;
wire [32*C_WIDTH-1:0] out_1419;
wire [32*C_WIDTH-1:0] out_1420;
wire [32*C_WIDTH-1:0] out_1421;
wire [32*C_WIDTH-1:0] out_1422;
wire [32*C_WIDTH-1:0] out_1423;
wire [32*C_WIDTH-1:0] out_1424;
wire [32*C_WIDTH-1:0] out_1425;
wire [32*C_WIDTH-1:0] out_1426;
wire [32*C_WIDTH-1:0] out_1427;
wire [32*C_WIDTH-1:0] out_1428;
wire [32*C_WIDTH-1:0] out_1429;
wire [32*C_WIDTH-1:0] out_1430;
wire [32*C_WIDTH-1:0] out_1431;
wire [32*C_WIDTH-1:0] out_1432;
wire [32*C_WIDTH-1:0] out_1433;
wire [32*C_WIDTH-1:0] out_1434;
wire [32*C_WIDTH-1:0] out_1435;
wire [32*C_WIDTH-1:0] out_1436;
wire [32*C_WIDTH-1:0] out_1437;
wire [32*C_WIDTH-1:0] out_1438;
wire [32*C_WIDTH-1:0] out_1439;
wire [32*C_WIDTH-1:0] out_1440;
wire [32*C_WIDTH-1:0] out_1441;
wire [32*C_WIDTH-1:0] out_1442;
wire [32*C_WIDTH-1:0] out_1443;
wire [32*C_WIDTH-1:0] out_1444;
wire [32*C_WIDTH-1:0] out_1445;
wire [32*C_WIDTH-1:0] out_1446;
wire [32*C_WIDTH-1:0] out_1447;
wire [32*C_WIDTH-1:0] out_1448;
wire [32*C_WIDTH-1:0] out_1449;
wire [32*C_WIDTH-1:0] out_1450;
wire [32*C_WIDTH-1:0] out_1451;
wire [32*C_WIDTH-1:0] out_1452;
wire [32*C_WIDTH-1:0] out_1453;
wire [32*C_WIDTH-1:0] out_1454;
wire [32*C_WIDTH-1:0] out_1455;
wire [32*C_WIDTH-1:0] out_1456;
wire [32*C_WIDTH-1:0] out_1457;
wire [32*C_WIDTH-1:0] out_1458;
wire [32*C_WIDTH-1:0] out_1459;
wire [32*C_WIDTH-1:0] out_1460;
wire [32*C_WIDTH-1:0] out_1461;
wire [32*C_WIDTH-1:0] out_1462;
wire [32*C_WIDTH-1:0] out_1463;
wire [32*C_WIDTH-1:0] out_1464;
wire [32*C_WIDTH-1:0] out_1465;
wire [32*C_WIDTH-1:0] out_1466;
wire [32*C_WIDTH-1:0] out_1467;
wire [32*C_WIDTH-1:0] out_1468;
wire [32*C_WIDTH-1:0] out_1469;
wire [32*C_WIDTH-1:0] out_1470;
wire [32*C_WIDTH-1:0] out_1471;
wire [32*C_WIDTH-1:0] out_1472;
wire [32*C_WIDTH-1:0] out_1473;
wire [32*C_WIDTH-1:0] out_1474;
wire [32*C_WIDTH-1:0] out_1475;
wire [32*C_WIDTH-1:0] out_1476;
wire [32*C_WIDTH-1:0] out_1477;
wire [32*C_WIDTH-1:0] out_1478;
wire [32*C_WIDTH-1:0] out_1479;
wire [32*C_WIDTH-1:0] out_1480;
wire [32*C_WIDTH-1:0] out_1481;
wire [32*C_WIDTH-1:0] out_1482;
wire [32*C_WIDTH-1:0] out_1483;
wire [32*C_WIDTH-1:0] out_1484;
wire [32*C_WIDTH-1:0] out_1485;
wire [32*C_WIDTH-1:0] out_1486;
wire [32*C_WIDTH-1:0] out_1487;
wire [32*C_WIDTH-1:0] out_1488;
wire [32*C_WIDTH-1:0] out_1489;
wire [32*C_WIDTH-1:0] out_1490;
wire [32*C_WIDTH-1:0] out_1491;
wire [32*C_WIDTH-1:0] out_1492;
wire [32*C_WIDTH-1:0] out_1493;
wire [32*C_WIDTH-1:0] out_1494;
wire [32*C_WIDTH-1:0] out_1495;
wire [32*C_WIDTH-1:0] out_1496;
wire [32*C_WIDTH-1:0] out_1497;
wire [32*C_WIDTH-1:0] out_1498;
wire [32*C_WIDTH-1:0] out_1499;
wire [32*C_WIDTH-1:0] out_1500;
wire [32*C_WIDTH-1:0] out_1501;
wire [32*C_WIDTH-1:0] out_1502;
wire [32*C_WIDTH-1:0] out_1503;
wire [32*C_WIDTH-1:0] out_1504;
wire [32*C_WIDTH-1:0] out_1505;
wire [32*C_WIDTH-1:0] out_1506;
wire [32*C_WIDTH-1:0] out_1507;
wire [32*C_WIDTH-1:0] out_1508;
wire [32*C_WIDTH-1:0] out_1509;
wire [32*C_WIDTH-1:0] out_1510;
wire [32*C_WIDTH-1:0] out_1511;
wire [32*C_WIDTH-1:0] out_1512;
wire [32*C_WIDTH-1:0] out_1513;
wire [32*C_WIDTH-1:0] out_1514;
wire [32*C_WIDTH-1:0] out_1515;
wire [32*C_WIDTH-1:0] out_1516;
wire [32*C_WIDTH-1:0] out_1517;
wire [32*C_WIDTH-1:0] out_1518;
wire [32*C_WIDTH-1:0] out_1519;
wire [32*C_WIDTH-1:0] out_1520;
wire [32*C_WIDTH-1:0] out_1521;
wire [32*C_WIDTH-1:0] out_1522;
wire [32*C_WIDTH-1:0] out_1523;
wire [32*C_WIDTH-1:0] out_1524;
wire [32*C_WIDTH-1:0] out_1525;
wire [32*C_WIDTH-1:0] out_1526;
wire [32*C_WIDTH-1:0] out_1527;
wire [32*C_WIDTH-1:0] out_1528;
wire [32*C_WIDTH-1:0] out_1529;
wire [32*C_WIDTH-1:0] out_1530;
wire [32*C_WIDTH-1:0] out_1531;
wire [32*C_WIDTH-1:0] out_1532;
wire [32*C_WIDTH-1:0] out_1533;
wire [32*C_WIDTH-1:0] out_1534;
wire [32*C_WIDTH-1:0] out_1535;
wire [32*C_WIDTH-1:0] out_1536;
wire [32*C_WIDTH-1:0] out_1537;
wire [32*C_WIDTH-1:0] out_1538;
wire [32*C_WIDTH-1:0] out_1539;
wire [32*C_WIDTH-1:0] out_1540;
wire [32*C_WIDTH-1:0] out_1541;
wire [32*C_WIDTH-1:0] out_1542;
wire [32*C_WIDTH-1:0] out_1543;
wire [32*C_WIDTH-1:0] out_1544;
wire [32*C_WIDTH-1:0] out_1545;
wire [32*C_WIDTH-1:0] out_1546;
wire [32*C_WIDTH-1:0] out_1547;
wire [32*C_WIDTH-1:0] out_1548;
wire [32*C_WIDTH-1:0] out_1549;
wire [32*C_WIDTH-1:0] out_1550;
wire [32*C_WIDTH-1:0] out_1551;
wire [32*C_WIDTH-1:0] out_1552;
wire [32*C_WIDTH-1:0] out_1553;
wire [32*C_WIDTH-1:0] out_1554;
wire [32*C_WIDTH-1:0] out_1555;
wire [32*C_WIDTH-1:0] out_1556;
wire [32*C_WIDTH-1:0] out_1557;
wire [32*C_WIDTH-1:0] out_1558;
wire [32*C_WIDTH-1:0] out_1559;
wire [32*C_WIDTH-1:0] out_1560;
wire [32*C_WIDTH-1:0] out_1561;
wire [32*C_WIDTH-1:0] out_1562;
wire [32*C_WIDTH-1:0] out_1563;
wire [32*C_WIDTH-1:0] out_1564;
wire [32*C_WIDTH-1:0] out_1565;
wire [32*C_WIDTH-1:0] out_1566;
wire [32*C_WIDTH-1:0] out_1567;
wire [32*C_WIDTH-1:0] out_1568;
wire [32*C_WIDTH-1:0] out_1569;
wire [32*C_WIDTH-1:0] out_1570;
wire [32*C_WIDTH-1:0] out_1571;
wire [32*C_WIDTH-1:0] out_1572;
wire [32*C_WIDTH-1:0] out_1573;
wire [32*C_WIDTH-1:0] out_1574;
wire [32*C_WIDTH-1:0] out_1575;
wire [32*C_WIDTH-1:0] out_1576;
wire [32*C_WIDTH-1:0] out_1577;
wire [32*C_WIDTH-1:0] out_1578;
wire [32*C_WIDTH-1:0] out_1579;
wire [32*C_WIDTH-1:0] out_1580;
wire [32*C_WIDTH-1:0] out_1581;
wire [32*C_WIDTH-1:0] out_1582;
wire [32*C_WIDTH-1:0] out_1583;
wire [32*C_WIDTH-1:0] out_1584;
wire [32*C_WIDTH-1:0] out_1585;
wire [32*C_WIDTH-1:0] out_1586;
wire [32*C_WIDTH-1:0] out_1587;
wire [32*C_WIDTH-1:0] out_1588;
wire [32*C_WIDTH-1:0] out_1589;
wire [32*C_WIDTH-1:0] out_1590;
wire [32*C_WIDTH-1:0] out_1591;
wire [32*C_WIDTH-1:0] out_1592;
wire [32*C_WIDTH-1:0] out_1593;
wire [32*C_WIDTH-1:0] out_1594;
wire [32*C_WIDTH-1:0] out_1595;
wire [32*C_WIDTH-1:0] out_1596;
wire [32*C_WIDTH-1:0] out_1597;
wire [32*C_WIDTH-1:0] out_1598;
wire [32*C_WIDTH-1:0] out_1599;
wire [32*C_WIDTH-1:0] out_1600;
wire [32*C_WIDTH-1:0] out_1601;
wire [32*C_WIDTH-1:0] out_1602;
wire [32*C_WIDTH-1:0] out_1603;
wire [32*C_WIDTH-1:0] out_1604;
wire [32*C_WIDTH-1:0] out_1605;
wire [32*C_WIDTH-1:0] out_1606;
wire [32*C_WIDTH-1:0] out_1607;
wire [32*C_WIDTH-1:0] out_1608;
wire [32*C_WIDTH-1:0] out_1609;
wire [32*C_WIDTH-1:0] out_1610;
wire [32*C_WIDTH-1:0] out_1611;
wire [32*C_WIDTH-1:0] out_1612;
wire [32*C_WIDTH-1:0] out_1613;
wire [32*C_WIDTH-1:0] out_1614;
wire [32*C_WIDTH-1:0] out_1615;
wire [32*C_WIDTH-1:0] out_1616;
wire [32*C_WIDTH-1:0] out_1617;
wire [32*C_WIDTH-1:0] out_1618;
wire [32*C_WIDTH-1:0] out_1619;
wire [32*C_WIDTH-1:0] out_1620;
wire [32*C_WIDTH-1:0] out_1621;
wire [32*C_WIDTH-1:0] out_1622;
wire [32*C_WIDTH-1:0] out_1623;
wire [32*C_WIDTH-1:0] out_1624;
wire [32*C_WIDTH-1:0] out_1625;
wire [32*C_WIDTH-1:0] out_1626;
wire [32*C_WIDTH-1:0] out_1627;
wire [32*C_WIDTH-1:0] out_1628;
wire [32*C_WIDTH-1:0] out_1629;
wire [32*C_WIDTH-1:0] out_1630;
wire [32*C_WIDTH-1:0] out_1631;
wire [32*C_WIDTH-1:0] out_1632;
wire [32*C_WIDTH-1:0] out_1633;
wire [32*C_WIDTH-1:0] out_1634;
wire [32*C_WIDTH-1:0] out_1635;
wire [32*C_WIDTH-1:0] out_1636;
wire [32*C_WIDTH-1:0] out_1637;
wire [32*C_WIDTH-1:0] out_1638;
wire [32*C_WIDTH-1:0] out_1639;
wire [32*C_WIDTH-1:0] out_1640;
wire [32*C_WIDTH-1:0] out_1641;
wire [32*C_WIDTH-1:0] out_1642;
wire [32*C_WIDTH-1:0] out_1643;
wire [32*C_WIDTH-1:0] out_1644;
wire [32*C_WIDTH-1:0] out_1645;
wire [32*C_WIDTH-1:0] out_1646;
wire [32*C_WIDTH-1:0] out_1647;
wire [32*C_WIDTH-1:0] out_1648;
wire [32*C_WIDTH-1:0] out_1649;
wire [32*C_WIDTH-1:0] out_1650;
wire [32*C_WIDTH-1:0] out_1651;
wire [32*C_WIDTH-1:0] out_1652;
wire [32*C_WIDTH-1:0] out_1653;
wire [32*C_WIDTH-1:0] out_1654;
wire [32*C_WIDTH-1:0] out_1655;
wire [32*C_WIDTH-1:0] out_1656;
wire [32*C_WIDTH-1:0] out_1657;
wire [32*C_WIDTH-1:0] out_1658;
wire [32*C_WIDTH-1:0] out_1659;
wire [32*C_WIDTH-1:0] out_1660;
wire [32*C_WIDTH-1:0] out_1661;
wire [32*C_WIDTH-1:0] out_1662;
wire [32*C_WIDTH-1:0] out_1663;
wire [32*C_WIDTH-1:0] out_1664;
wire [32*C_WIDTH-1:0] out_1665;
wire [32*C_WIDTH-1:0] out_1666;
wire [32*C_WIDTH-1:0] out_1667;
wire [32*C_WIDTH-1:0] out_1668;
wire [32*C_WIDTH-1:0] out_1669;
wire [32*C_WIDTH-1:0] out_1670;
wire [32*C_WIDTH-1:0] out_1671;
wire [32*C_WIDTH-1:0] out_1672;
wire [32*C_WIDTH-1:0] out_1673;
wire [32*C_WIDTH-1:0] out_1674;
wire [32*C_WIDTH-1:0] out_1675;
wire [32*C_WIDTH-1:0] out_1676;
wire [32*C_WIDTH-1:0] out_1677;
wire [32*C_WIDTH-1:0] out_1678;
wire [32*C_WIDTH-1:0] out_1679;
wire [32*C_WIDTH-1:0] out_1680;
wire [32*C_WIDTH-1:0] out_1681;
wire [32*C_WIDTH-1:0] out_1682;
wire [32*C_WIDTH-1:0] out_1683;
wire [32*C_WIDTH-1:0] out_1684;
wire [32*C_WIDTH-1:0] out_1685;
wire [32*C_WIDTH-1:0] out_1686;
wire [32*C_WIDTH-1:0] out_1687;
wire [32*C_WIDTH-1:0] out_1688;
wire [32*C_WIDTH-1:0] out_1689;
wire [32*C_WIDTH-1:0] out_1690;
wire [32*C_WIDTH-1:0] out_1691;
wire [32*C_WIDTH-1:0] out_1692;
wire [32*C_WIDTH-1:0] out_1693;
wire [32*C_WIDTH-1:0] out_1694;
wire [32*C_WIDTH-1:0] out_1695;
wire [32*C_WIDTH-1:0] out_1696;
wire [32*C_WIDTH-1:0] out_1697;
wire [32*C_WIDTH-1:0] out_1698;
wire [32*C_WIDTH-1:0] out_1699;
wire [32*C_WIDTH-1:0] out_1700;
wire [32*C_WIDTH-1:0] out_1701;
wire [32*C_WIDTH-1:0] out_1702;
wire [32*C_WIDTH-1:0] out_1703;
wire [32*C_WIDTH-1:0] out_1704;
wire [32*C_WIDTH-1:0] out_1705;
wire [32*C_WIDTH-1:0] out_1706;
wire [32*C_WIDTH-1:0] out_1707;
wire [32*C_WIDTH-1:0] out_1708;
wire [32*C_WIDTH-1:0] out_1709;
wire [32*C_WIDTH-1:0] out_1710;
wire [32*C_WIDTH-1:0] out_1711;
wire [32*C_WIDTH-1:0] out_1712;
wire [32*C_WIDTH-1:0] out_1713;
wire [32*C_WIDTH-1:0] out_1714;
wire [32*C_WIDTH-1:0] out_1715;
wire [32*C_WIDTH-1:0] out_1716;
wire [32*C_WIDTH-1:0] out_1717;
wire [32*C_WIDTH-1:0] out_1718;
wire [32*C_WIDTH-1:0] out_1719;
wire [32*C_WIDTH-1:0] out_1720;
wire [32*C_WIDTH-1:0] out_1721;
wire [32*C_WIDTH-1:0] out_1722;
wire [32*C_WIDTH-1:0] out_1723;
wire [32*C_WIDTH-1:0] out_1724;
wire [32*C_WIDTH-1:0] out_1725;
wire [32*C_WIDTH-1:0] out_1726;
wire [32*C_WIDTH-1:0] out_1727;
wire [32*C_WIDTH-1:0] out_1728;
wire [32*C_WIDTH-1:0] out_1729;
wire [32*C_WIDTH-1:0] out_1730;
wire [32*C_WIDTH-1:0] out_1731;
wire [32*C_WIDTH-1:0] out_1732;
wire [32*C_WIDTH-1:0] out_1733;
wire [32*C_WIDTH-1:0] out_1734;
wire [32*C_WIDTH-1:0] out_1735;
wire [32*C_WIDTH-1:0] out_1736;
wire [32*C_WIDTH-1:0] out_1737;
wire [32*C_WIDTH-1:0] out_1738;
wire [32*C_WIDTH-1:0] out_1739;
wire [32*C_WIDTH-1:0] out_1740;
wire [32*C_WIDTH-1:0] out_1741;
wire [32*C_WIDTH-1:0] out_1742;
wire [32*C_WIDTH-1:0] out_1743;
wire [32*C_WIDTH-1:0] out_1744;
wire [32*C_WIDTH-1:0] out_1745;
wire [32*C_WIDTH-1:0] out_1746;
wire [32*C_WIDTH-1:0] out_1747;
wire [32*C_WIDTH-1:0] out_1748;
wire [32*C_WIDTH-1:0] out_1749;
wire [32*C_WIDTH-1:0] out_1750;
wire [32*C_WIDTH-1:0] out_1751;
wire [32*C_WIDTH-1:0] out_1752;
wire [32*C_WIDTH-1:0] out_1753;
wire [32*C_WIDTH-1:0] out_1754;
wire [32*C_WIDTH-1:0] out_1755;
wire [32*C_WIDTH-1:0] out_1756;
wire [32*C_WIDTH-1:0] out_1757;
wire [32*C_WIDTH-1:0] out_1758;
wire [32*C_WIDTH-1:0] out_1759;
wire [32*C_WIDTH-1:0] out_1760;
wire [32*C_WIDTH-1:0] out_1761;
wire [32*C_WIDTH-1:0] out_1762;
wire [32*C_WIDTH-1:0] out_1763;
wire [32*C_WIDTH-1:0] out_1764;
wire [32*C_WIDTH-1:0] out_1765;
wire [32*C_WIDTH-1:0] out_1766;
wire [32*C_WIDTH-1:0] out_1767;
wire [32*C_WIDTH-1:0] out_1768;
wire [32*C_WIDTH-1:0] out_1769;
wire [32*C_WIDTH-1:0] out_1770;
wire [32*C_WIDTH-1:0] out_1771;
wire [32*C_WIDTH-1:0] out_1772;
wire [32*C_WIDTH-1:0] out_1773;
wire [32*C_WIDTH-1:0] out_1774;
wire [32*C_WIDTH-1:0] out_1775;
wire [32*C_WIDTH-1:0] out_1776;
wire [32*C_WIDTH-1:0] out_1777;
wire [32*C_WIDTH-1:0] out_1778;
wire [32*C_WIDTH-1:0] out_1779;
wire [32*C_WIDTH-1:0] out_1780;
wire [32*C_WIDTH-1:0] out_1781;
wire [32*C_WIDTH-1:0] out_1782;
wire [32*C_WIDTH-1:0] out_1783;
wire [32*C_WIDTH-1:0] out_1784;
wire [32*C_WIDTH-1:0] out_1785;
wire [32*C_WIDTH-1:0] out_1786;
wire [32*C_WIDTH-1:0] out_1787;
wire [32*C_WIDTH-1:0] out_1788;
wire [32*C_WIDTH-1:0] out_1789;
wire [32*C_WIDTH-1:0] out_1790;
wire [32*C_WIDTH-1:0] out_1791;
wire [32*C_WIDTH-1:0] out_1792;
wire [32*C_WIDTH-1:0] out_1793;
wire [32*C_WIDTH-1:0] out_1794;
wire [32*C_WIDTH-1:0] out_1795;
wire [32*C_WIDTH-1:0] out_1796;
wire [32*C_WIDTH-1:0] out_1797;
wire [32*C_WIDTH-1:0] out_1798;
wire [32*C_WIDTH-1:0] out_1799;
wire [32*C_WIDTH-1:0] out_1800;
wire [32*C_WIDTH-1:0] out_1801;
wire [32*C_WIDTH-1:0] out_1802;
wire [32*C_WIDTH-1:0] out_1803;
wire [32*C_WIDTH-1:0] out_1804;
wire [32*C_WIDTH-1:0] out_1805;
wire [32*C_WIDTH-1:0] out_1806;
wire [32*C_WIDTH-1:0] out_1807;
wire [32*C_WIDTH-1:0] out_1808;
wire [32*C_WIDTH-1:0] out_1809;
wire [32*C_WIDTH-1:0] out_1810;
wire [32*C_WIDTH-1:0] out_1811;
wire [32*C_WIDTH-1:0] out_1812;
wire [32*C_WIDTH-1:0] out_1813;
wire [32*C_WIDTH-1:0] out_1814;
wire [32*C_WIDTH-1:0] out_1815;
wire [32*C_WIDTH-1:0] out_1816;
wire [32*C_WIDTH-1:0] out_1817;
wire [32*C_WIDTH-1:0] out_1818;
wire [32*C_WIDTH-1:0] out_1819;
wire [32*C_WIDTH-1:0] out_1820;
wire [32*C_WIDTH-1:0] out_1821;
wire [32*C_WIDTH-1:0] out_1822;
wire [32*C_WIDTH-1:0] out_1823;
wire [32*C_WIDTH-1:0] out_1824;
wire [32*C_WIDTH-1:0] out_1825;
wire [32*C_WIDTH-1:0] out_1826;
wire [32*C_WIDTH-1:0] out_1827;
wire [32*C_WIDTH-1:0] out_1828;
wire [32*C_WIDTH-1:0] out_1829;
wire [32*C_WIDTH-1:0] out_1830;
wire [32*C_WIDTH-1:0] out_1831;
wire [32*C_WIDTH-1:0] out_1832;
wire [32*C_WIDTH-1:0] out_1833;
wire [32*C_WIDTH-1:0] out_1834;
wire [32*C_WIDTH-1:0] out_1835;
wire [32*C_WIDTH-1:0] out_1836;
wire [32*C_WIDTH-1:0] out_1837;
wire [32*C_WIDTH-1:0] out_1838;
wire [32*C_WIDTH-1:0] out_1839;
wire [32*C_WIDTH-1:0] out_1840;
wire [32*C_WIDTH-1:0] out_1841;
wire [32*C_WIDTH-1:0] out_1842;
wire [32*C_WIDTH-1:0] out_1843;
wire [32*C_WIDTH-1:0] out_1844;
wire [32*C_WIDTH-1:0] out_1845;
wire [32*C_WIDTH-1:0] out_1846;
wire [32*C_WIDTH-1:0] out_1847;
wire [32*C_WIDTH-1:0] out_1848;
wire [32*C_WIDTH-1:0] out_1849;
wire [32*C_WIDTH-1:0] out_1850;
wire [32*C_WIDTH-1:0] out_1851;
wire [32*C_WIDTH-1:0] out_1852;
wire [32*C_WIDTH-1:0] out_1853;
wire [32*C_WIDTH-1:0] out_1854;
wire [32*C_WIDTH-1:0] out_1855;
wire [32*C_WIDTH-1:0] out_1856;
wire [32*C_WIDTH-1:0] out_1857;
wire [32*C_WIDTH-1:0] out_1858;
wire [32*C_WIDTH-1:0] out_1859;
wire [32*C_WIDTH-1:0] out_1860;
wire [32*C_WIDTH-1:0] out_1861;
wire [32*C_WIDTH-1:0] out_1862;
wire [32*C_WIDTH-1:0] out_1863;
wire [32*C_WIDTH-1:0] out_1864;
wire [32*C_WIDTH-1:0] out_1865;
wire [32*C_WIDTH-1:0] out_1866;
wire [32*C_WIDTH-1:0] out_1867;
wire [32*C_WIDTH-1:0] out_1868;
wire [32*C_WIDTH-1:0] out_1869;
wire [32*C_WIDTH-1:0] out_1870;
wire [32*C_WIDTH-1:0] out_1871;
wire [32*C_WIDTH-1:0] out_1872;
wire [32*C_WIDTH-1:0] out_1873;
wire [32*C_WIDTH-1:0] out_1874;
wire [32*C_WIDTH-1:0] out_1875;
wire [32*C_WIDTH-1:0] out_1876;
wire [32*C_WIDTH-1:0] out_1877;
wire [32*C_WIDTH-1:0] out_1878;
wire [32*C_WIDTH-1:0] out_1879;
wire [32*C_WIDTH-1:0] out_1880;
wire [32*C_WIDTH-1:0] out_1881;
wire [32*C_WIDTH-1:0] out_1882;
wire [32*C_WIDTH-1:0] out_1883;
wire [32*C_WIDTH-1:0] out_1884;
wire [32*C_WIDTH-1:0] out_1885;
wire [32*C_WIDTH-1:0] out_1886;
wire [32*C_WIDTH-1:0] out_1887;
wire [32*C_WIDTH-1:0] out_1888;
wire [32*C_WIDTH-1:0] out_1889;
wire [32*C_WIDTH-1:0] out_1890;
wire [32*C_WIDTH-1:0] out_1891;
wire [32*C_WIDTH-1:0] out_1892;
wire [32*C_WIDTH-1:0] out_1893;
wire [32*C_WIDTH-1:0] out_1894;
wire [32*C_WIDTH-1:0] out_1895;
wire [32*C_WIDTH-1:0] out_1896;
wire [32*C_WIDTH-1:0] out_1897;
wire [32*C_WIDTH-1:0] out_1898;
wire [32*C_WIDTH-1:0] out_1899;
wire [32*C_WIDTH-1:0] out_1900;
wire [32*C_WIDTH-1:0] out_1901;
wire [32*C_WIDTH-1:0] out_1902;
wire [32*C_WIDTH-1:0] out_1903;
wire [32*C_WIDTH-1:0] out_1904;
wire [32*C_WIDTH-1:0] out_1905;
wire [32*C_WIDTH-1:0] out_1906;
wire [32*C_WIDTH-1:0] out_1907;
wire [32*C_WIDTH-1:0] out_1908;
wire [32*C_WIDTH-1:0] out_1909;
wire [32*C_WIDTH-1:0] out_1910;
wire [32*C_WIDTH-1:0] out_1911;
wire [32*C_WIDTH-1:0] out_1912;
wire [32*C_WIDTH-1:0] out_1913;
wire [32*C_WIDTH-1:0] out_1914;
wire [32*C_WIDTH-1:0] out_1915;
wire [32*C_WIDTH-1:0] out_1916;
wire [32*C_WIDTH-1:0] out_1917;
wire [32*C_WIDTH-1:0] out_1918;
wire [32*C_WIDTH-1:0] out_1919;
wire [32*C_WIDTH-1:0] out_1920;
wire [32*C_WIDTH-1:0] out_1921;
wire [32*C_WIDTH-1:0] out_1922;
wire [32*C_WIDTH-1:0] out_1923;
wire [32*C_WIDTH-1:0] out_1924;
wire [32*C_WIDTH-1:0] out_1925;
wire [32*C_WIDTH-1:0] out_1926;
wire [32*C_WIDTH-1:0] out_1927;
wire [32*C_WIDTH-1:0] out_1928;
wire [32*C_WIDTH-1:0] out_1929;
wire [32*C_WIDTH-1:0] out_1930;
wire [32*C_WIDTH-1:0] out_1931;
wire [32*C_WIDTH-1:0] out_1932;
wire [32*C_WIDTH-1:0] out_1933;
wire [32*C_WIDTH-1:0] out_1934;
wire [32*C_WIDTH-1:0] out_1935;
wire [32*C_WIDTH-1:0] out_1936;
wire [32*C_WIDTH-1:0] out_1937;
wire [32*C_WIDTH-1:0] out_1938;
wire [32*C_WIDTH-1:0] out_1939;
wire [32*C_WIDTH-1:0] out_1940;
wire [32*C_WIDTH-1:0] out_1941;
wire [32*C_WIDTH-1:0] out_1942;
wire [32*C_WIDTH-1:0] out_1943;
wire [32*C_WIDTH-1:0] out_1944;
wire [32*C_WIDTH-1:0] out_1945;
wire [32*C_WIDTH-1:0] out_1946;
wire [32*C_WIDTH-1:0] out_1947;
wire [32*C_WIDTH-1:0] out_1948;
wire [32*C_WIDTH-1:0] out_1949;
wire [32*C_WIDTH-1:0] out_1950;
wire [32*C_WIDTH-1:0] out_1951;
wire [32*C_WIDTH-1:0] out_1952;
wire [32*C_WIDTH-1:0] out_1953;
wire [32*C_WIDTH-1:0] out_1954;
wire [32*C_WIDTH-1:0] out_1955;
wire [32*C_WIDTH-1:0] out_1956;
wire [32*C_WIDTH-1:0] out_1957;
wire [32*C_WIDTH-1:0] out_1958;
wire [32*C_WIDTH-1:0] out_1959;
wire [32*C_WIDTH-1:0] out_1960;
wire [32*C_WIDTH-1:0] out_1961;
wire [32*C_WIDTH-1:0] out_1962;
wire [32*C_WIDTH-1:0] out_1963;
wire [32*C_WIDTH-1:0] out_1964;
wire [32*C_WIDTH-1:0] out_1965;
wire [32*C_WIDTH-1:0] out_1966;
wire [32*C_WIDTH-1:0] out_1967;
wire [32*C_WIDTH-1:0] out_1968;
wire [32*C_WIDTH-1:0] out_1969;
wire [32*C_WIDTH-1:0] out_1970;
wire [32*C_WIDTH-1:0] out_1971;
wire [32*C_WIDTH-1:0] out_1972;
wire [32*C_WIDTH-1:0] out_1973;
wire [32*C_WIDTH-1:0] out_1974;
wire [32*C_WIDTH-1:0] out_1975;
wire [32*C_WIDTH-1:0] out_1976;
wire [32*C_WIDTH-1:0] out_1977;
wire [32*C_WIDTH-1:0] out_1978;
wire [32*C_WIDTH-1:0] out_1979;
wire [32*C_WIDTH-1:0] out_1980;
wire [32*C_WIDTH-1:0] out_1981;
wire [32*C_WIDTH-1:0] out_1982;
wire [32*C_WIDTH-1:0] out_1983;
wire [32*C_WIDTH-1:0] out_1984;
wire [32*C_WIDTH-1:0] out_1985;
wire [32*C_WIDTH-1:0] out_1986;
wire [32*C_WIDTH-1:0] out_1987;
wire [32*C_WIDTH-1:0] out_1988;
wire [32*C_WIDTH-1:0] out_1989;
wire [32*C_WIDTH-1:0] out_1990;
wire [32*C_WIDTH-1:0] out_1991;
wire [32*C_WIDTH-1:0] out_1992;
wire [32*C_WIDTH-1:0] out_1993;
wire [32*C_WIDTH-1:0] out_1994;
wire [32*C_WIDTH-1:0] out_1995;
wire [32*C_WIDTH-1:0] out_1996;
wire [32*C_WIDTH-1:0] out_1997;
wire [32*C_WIDTH-1:0] out_1998;
wire [32*C_WIDTH-1:0] out_1999;
wire [32*C_WIDTH-1:0] out_2000;
wire [32*C_WIDTH-1:0] out_2001;
wire [32*C_WIDTH-1:0] out_2002;
wire [32*C_WIDTH-1:0] out_2003;
wire [32*C_WIDTH-1:0] out_2004;
wire [32*C_WIDTH-1:0] out_2005;
wire [32*C_WIDTH-1:0] out_2006;
wire [32*C_WIDTH-1:0] out_2007;
wire [32*C_WIDTH-1:0] out_2008;
wire [32*C_WIDTH-1:0] out_2009;
wire [32*C_WIDTH-1:0] out_2010;
wire [32*C_WIDTH-1:0] out_2011;
wire [32*C_WIDTH-1:0] out_2012;
wire [32*C_WIDTH-1:0] out_2013;
wire [32*C_WIDTH-1:0] out_2014;
wire [32*C_WIDTH-1:0] out_2015;
wire [32*C_WIDTH-1:0] out_2016;
wire [32*C_WIDTH-1:0] out_2017;
wire [32*C_WIDTH-1:0] out_2018;
wire [32*C_WIDTH-1:0] out_2019;
wire [32*C_WIDTH-1:0] out_2020;
wire [32*C_WIDTH-1:0] out_2021;
wire [32*C_WIDTH-1:0] out_2022;
wire [32*C_WIDTH-1:0] out_2023;
wire [32*C_WIDTH-1:0] out_2024;
wire [32*C_WIDTH-1:0] out_2025;
wire [32*C_WIDTH-1:0] out_2026;
wire [32*C_WIDTH-1:0] out_2027;
wire [32*C_WIDTH-1:0] out_2028;
wire [32*C_WIDTH-1:0] out_2029;
wire [32*C_WIDTH-1:0] out_2030;
wire [32*C_WIDTH-1:0] out_2031;
wire [32*C_WIDTH-1:0] out_2032;
wire [32*C_WIDTH-1:0] out_2033;
wire [32*C_WIDTH-1:0] out_2034;
wire [32*C_WIDTH-1:0] out_2035;
wire [32*C_WIDTH-1:0] out_2036;
wire [32*C_WIDTH-1:0] out_2037;
wire [32*C_WIDTH-1:0] out_2038;
wire [32*C_WIDTH-1:0] out_2039;
wire [32*C_WIDTH-1:0] out_2040;
wire [32*C_WIDTH-1:0] out_2041;
wire [32*C_WIDTH-1:0] out_2042;
wire [32*C_WIDTH-1:0] out_2043;
wire [32*C_WIDTH-1:0] out_2044;
wire [32*C_WIDTH-1:0] out_2045;
wire [32*C_WIDTH-1:0] out_2046;
wire [32*C_WIDTH-1:0] out_2047;
assign {act_0,act_1} = activation;
assign {weight_0,weight_1} = weight;

SA128 SA128_0 (.clk(clk),.rstn(rstn),.activation(act_0),.weight(weight_0),.out_act(act0_1),.out_weight(weight0_2),.control(control),.c_out0(out_0),
.c_out1(out_1),
.c_out2(out_2),
.c_out3(out_3),
.c_out4(out_4),
.c_out5(out_5),
.c_out6(out_6),
.c_out7(out_7),
.c_out8(out_8),
.c_out9(out_9),
.c_out10(out_10),
.c_out11(out_11),
.c_out12(out_12),
.c_out13(out_13),
.c_out14(out_14),
.c_out15(out_15),
.c_out16(out_16),
.c_out17(out_17),
.c_out18(out_18),
.c_out19(out_19),
.c_out20(out_20),
.c_out21(out_21),
.c_out22(out_22),
.c_out23(out_23),
.c_out24(out_24),
.c_out25(out_25),
.c_out26(out_26),
.c_out27(out_27),
.c_out28(out_28),
.c_out29(out_29),
.c_out30(out_30),
.c_out31(out_31),
.c_out32(out_32),
.c_out33(out_33),
.c_out34(out_34),
.c_out35(out_35),
.c_out36(out_36),
.c_out37(out_37),
.c_out38(out_38),
.c_out39(out_39),
.c_out40(out_40),
.c_out41(out_41),
.c_out42(out_42),
.c_out43(out_43),
.c_out44(out_44),
.c_out45(out_45),
.c_out46(out_46),
.c_out47(out_47),
.c_out48(out_48),
.c_out49(out_49),
.c_out50(out_50),
.c_out51(out_51),
.c_out52(out_52),
.c_out53(out_53),
.c_out54(out_54),
.c_out55(out_55),
.c_out56(out_56),
.c_out57(out_57),
.c_out58(out_58),
.c_out59(out_59),
.c_out60(out_60),
.c_out61(out_61),
.c_out62(out_62),
.c_out63(out_63),
.c_out64(out_64),
.c_out65(out_65),
.c_out66(out_66),
.c_out67(out_67),
.c_out68(out_68),
.c_out69(out_69),
.c_out70(out_70),
.c_out71(out_71),
.c_out72(out_72),
.c_out73(out_73),
.c_out74(out_74),
.c_out75(out_75),
.c_out76(out_76),
.c_out77(out_77),
.c_out78(out_78),
.c_out79(out_79),
.c_out80(out_80),
.c_out81(out_81),
.c_out82(out_82),
.c_out83(out_83),
.c_out84(out_84),
.c_out85(out_85),
.c_out86(out_86),
.c_out87(out_87),
.c_out88(out_88),
.c_out89(out_89),
.c_out90(out_90),
.c_out91(out_91),
.c_out92(out_92),
.c_out93(out_93),
.c_out94(out_94),
.c_out95(out_95),
.c_out96(out_96),
.c_out97(out_97),
.c_out98(out_98),
.c_out99(out_99),
.c_out100(out_100),
.c_out101(out_101),
.c_out102(out_102),
.c_out103(out_103),
.c_out104(out_104),
.c_out105(out_105),
.c_out106(out_106),
.c_out107(out_107),
.c_out108(out_108),
.c_out109(out_109),
.c_out110(out_110),
.c_out111(out_111),
.c_out112(out_112),
.c_out113(out_113),
.c_out114(out_114),
.c_out115(out_115),
.c_out116(out_116),
.c_out117(out_117),
.c_out118(out_118),
.c_out119(out_119),
.c_out120(out_120),
.c_out121(out_121),
.c_out122(out_122),
.c_out123(out_123),
.c_out124(out_124),
.c_out125(out_125),
.c_out126(out_126),
.c_out127(out_127),
.c_out128(out_128),
.c_out129(out_129),
.c_out130(out_130),
.c_out131(out_131),
.c_out132(out_132),
.c_out133(out_133),
.c_out134(out_134),
.c_out135(out_135),
.c_out136(out_136),
.c_out137(out_137),
.c_out138(out_138),
.c_out139(out_139),
.c_out140(out_140),
.c_out141(out_141),
.c_out142(out_142),
.c_out143(out_143),
.c_out144(out_144),
.c_out145(out_145),
.c_out146(out_146),
.c_out147(out_147),
.c_out148(out_148),
.c_out149(out_149),
.c_out150(out_150),
.c_out151(out_151),
.c_out152(out_152),
.c_out153(out_153),
.c_out154(out_154),
.c_out155(out_155),
.c_out156(out_156),
.c_out157(out_157),
.c_out158(out_158),
.c_out159(out_159),
.c_out160(out_160),
.c_out161(out_161),
.c_out162(out_162),
.c_out163(out_163),
.c_out164(out_164),
.c_out165(out_165),
.c_out166(out_166),
.c_out167(out_167),
.c_out168(out_168),
.c_out169(out_169),
.c_out170(out_170),
.c_out171(out_171),
.c_out172(out_172),
.c_out173(out_173),
.c_out174(out_174),
.c_out175(out_175),
.c_out176(out_176),
.c_out177(out_177),
.c_out178(out_178),
.c_out179(out_179),
.c_out180(out_180),
.c_out181(out_181),
.c_out182(out_182),
.c_out183(out_183),
.c_out184(out_184),
.c_out185(out_185),
.c_out186(out_186),
.c_out187(out_187),
.c_out188(out_188),
.c_out189(out_189),
.c_out190(out_190),
.c_out191(out_191),
.c_out192(out_192),
.c_out193(out_193),
.c_out194(out_194),
.c_out195(out_195),
.c_out196(out_196),
.c_out197(out_197),
.c_out198(out_198),
.c_out199(out_199),
.c_out200(out_200),
.c_out201(out_201),
.c_out202(out_202),
.c_out203(out_203),
.c_out204(out_204),
.c_out205(out_205),
.c_out206(out_206),
.c_out207(out_207),
.c_out208(out_208),
.c_out209(out_209),
.c_out210(out_210),
.c_out211(out_211),
.c_out212(out_212),
.c_out213(out_213),
.c_out214(out_214),
.c_out215(out_215),
.c_out216(out_216),
.c_out217(out_217),
.c_out218(out_218),
.c_out219(out_219),
.c_out220(out_220),
.c_out221(out_221),
.c_out222(out_222),
.c_out223(out_223),
.c_out224(out_224),
.c_out225(out_225),
.c_out226(out_226),
.c_out227(out_227),
.c_out228(out_228),
.c_out229(out_229),
.c_out230(out_230),
.c_out231(out_231),
.c_out232(out_232),
.c_out233(out_233),
.c_out234(out_234),
.c_out235(out_235),
.c_out236(out_236),
.c_out237(out_237),
.c_out238(out_238),
.c_out239(out_239),
.c_out240(out_240),
.c_out241(out_241),
.c_out242(out_242),
.c_out243(out_243),
.c_out244(out_244),
.c_out245(out_245),
.c_out246(out_246),
.c_out247(out_247),
.c_out248(out_248),
.c_out249(out_249),
.c_out250(out_250),
.c_out251(out_251),
.c_out252(out_252),
.c_out253(out_253),
.c_out254(out_254),
.c_out255(out_255),
.c_out256(out_256),
.c_out257(out_257),
.c_out258(out_258),
.c_out259(out_259),
.c_out260(out_260),
.c_out261(out_261),
.c_out262(out_262),
.c_out263(out_263),
.c_out264(out_264),
.c_out265(out_265),
.c_out266(out_266),
.c_out267(out_267),
.c_out268(out_268),
.c_out269(out_269),
.c_out270(out_270),
.c_out271(out_271),
.c_out272(out_272),
.c_out273(out_273),
.c_out274(out_274),
.c_out275(out_275),
.c_out276(out_276),
.c_out277(out_277),
.c_out278(out_278),
.c_out279(out_279),
.c_out280(out_280),
.c_out281(out_281),
.c_out282(out_282),
.c_out283(out_283),
.c_out284(out_284),
.c_out285(out_285),
.c_out286(out_286),
.c_out287(out_287),
.c_out288(out_288),
.c_out289(out_289),
.c_out290(out_290),
.c_out291(out_291),
.c_out292(out_292),
.c_out293(out_293),
.c_out294(out_294),
.c_out295(out_295),
.c_out296(out_296),
.c_out297(out_297),
.c_out298(out_298),
.c_out299(out_299),
.c_out300(out_300),
.c_out301(out_301),
.c_out302(out_302),
.c_out303(out_303),
.c_out304(out_304),
.c_out305(out_305),
.c_out306(out_306),
.c_out307(out_307),
.c_out308(out_308),
.c_out309(out_309),
.c_out310(out_310),
.c_out311(out_311),
.c_out312(out_312),
.c_out313(out_313),
.c_out314(out_314),
.c_out315(out_315),
.c_out316(out_316),
.c_out317(out_317),
.c_out318(out_318),
.c_out319(out_319),
.c_out320(out_320),
.c_out321(out_321),
.c_out322(out_322),
.c_out323(out_323),
.c_out324(out_324),
.c_out325(out_325),
.c_out326(out_326),
.c_out327(out_327),
.c_out328(out_328),
.c_out329(out_329),
.c_out330(out_330),
.c_out331(out_331),
.c_out332(out_332),
.c_out333(out_333),
.c_out334(out_334),
.c_out335(out_335),
.c_out336(out_336),
.c_out337(out_337),
.c_out338(out_338),
.c_out339(out_339),
.c_out340(out_340),
.c_out341(out_341),
.c_out342(out_342),
.c_out343(out_343),
.c_out344(out_344),
.c_out345(out_345),
.c_out346(out_346),
.c_out347(out_347),
.c_out348(out_348),
.c_out349(out_349),
.c_out350(out_350),
.c_out351(out_351),
.c_out352(out_352),
.c_out353(out_353),
.c_out354(out_354),
.c_out355(out_355),
.c_out356(out_356),
.c_out357(out_357),
.c_out358(out_358),
.c_out359(out_359),
.c_out360(out_360),
.c_out361(out_361),
.c_out362(out_362),
.c_out363(out_363),
.c_out364(out_364),
.c_out365(out_365),
.c_out366(out_366),
.c_out367(out_367),
.c_out368(out_368),
.c_out369(out_369),
.c_out370(out_370),
.c_out371(out_371),
.c_out372(out_372),
.c_out373(out_373),
.c_out374(out_374),
.c_out375(out_375),
.c_out376(out_376),
.c_out377(out_377),
.c_out378(out_378),
.c_out379(out_379),
.c_out380(out_380),
.c_out381(out_381),
.c_out382(out_382),
.c_out383(out_383),
.c_out384(out_384),
.c_out385(out_385),
.c_out386(out_386),
.c_out387(out_387),
.c_out388(out_388),
.c_out389(out_389),
.c_out390(out_390),
.c_out391(out_391),
.c_out392(out_392),
.c_out393(out_393),
.c_out394(out_394),
.c_out395(out_395),
.c_out396(out_396),
.c_out397(out_397),
.c_out398(out_398),
.c_out399(out_399),
.c_out400(out_400),
.c_out401(out_401),
.c_out402(out_402),
.c_out403(out_403),
.c_out404(out_404),
.c_out405(out_405),
.c_out406(out_406),
.c_out407(out_407),
.c_out408(out_408),
.c_out409(out_409),
.c_out410(out_410),
.c_out411(out_411),
.c_out412(out_412),
.c_out413(out_413),
.c_out414(out_414),
.c_out415(out_415),
.c_out416(out_416),
.c_out417(out_417),
.c_out418(out_418),
.c_out419(out_419),
.c_out420(out_420),
.c_out421(out_421),
.c_out422(out_422),
.c_out423(out_423),
.c_out424(out_424),
.c_out425(out_425),
.c_out426(out_426),
.c_out427(out_427),
.c_out428(out_428),
.c_out429(out_429),
.c_out430(out_430),
.c_out431(out_431),
.c_out432(out_432),
.c_out433(out_433),
.c_out434(out_434),
.c_out435(out_435),
.c_out436(out_436),
.c_out437(out_437),
.c_out438(out_438),
.c_out439(out_439),
.c_out440(out_440),
.c_out441(out_441),
.c_out442(out_442),
.c_out443(out_443),
.c_out444(out_444),
.c_out445(out_445),
.c_out446(out_446),
.c_out447(out_447),
.c_out448(out_448),
.c_out449(out_449),
.c_out450(out_450),
.c_out451(out_451),
.c_out452(out_452),
.c_out453(out_453),
.c_out454(out_454),
.c_out455(out_455),
.c_out456(out_456),
.c_out457(out_457),
.c_out458(out_458),
.c_out459(out_459),
.c_out460(out_460),
.c_out461(out_461),
.c_out462(out_462),
.c_out463(out_463),
.c_out464(out_464),
.c_out465(out_465),
.c_out466(out_466),
.c_out467(out_467),
.c_out468(out_468),
.c_out469(out_469),
.c_out470(out_470),
.c_out471(out_471),
.c_out472(out_472),
.c_out473(out_473),
.c_out474(out_474),
.c_out475(out_475),
.c_out476(out_476),
.c_out477(out_477),
.c_out478(out_478),
.c_out479(out_479),
.c_out480(out_480),
.c_out481(out_481),
.c_out482(out_482),
.c_out483(out_483),
.c_out484(out_484),
.c_out485(out_485),
.c_out486(out_486),
.c_out487(out_487),
.c_out488(out_488),
.c_out489(out_489),
.c_out490(out_490),
.c_out491(out_491),
.c_out492(out_492),
.c_out493(out_493),
.c_out494(out_494),
.c_out495(out_495),
.c_out496(out_496),
.c_out497(out_497),
.c_out498(out_498),
.c_out499(out_499),
.c_out500(out_500),
.c_out501(out_501),
.c_out502(out_502),
.c_out503(out_503),
.c_out504(out_504),
.c_out505(out_505),
.c_out506(out_506),
.c_out507(out_507),
.c_out508(out_508),
.c_out509(out_509),
.c_out510(out_510),
.c_out511(out_511));
SA128 SA128_1 (.clk(clk),.rstn(rstn),.activation(act0_1),.weight(weight_1),.out_act(outact_0),.out_weight(weight1_3),.control(control),.c_out0(out_512),
.c_out1(out_513),
.c_out2(out_514),
.c_out3(out_515),
.c_out4(out_516),
.c_out5(out_517),
.c_out6(out_518),
.c_out7(out_519),
.c_out8(out_520),
.c_out9(out_521),
.c_out10(out_522),
.c_out11(out_523),
.c_out12(out_524),
.c_out13(out_525),
.c_out14(out_526),
.c_out15(out_527),
.c_out16(out_528),
.c_out17(out_529),
.c_out18(out_530),
.c_out19(out_531),
.c_out20(out_532),
.c_out21(out_533),
.c_out22(out_534),
.c_out23(out_535),
.c_out24(out_536),
.c_out25(out_537),
.c_out26(out_538),
.c_out27(out_539),
.c_out28(out_540),
.c_out29(out_541),
.c_out30(out_542),
.c_out31(out_543),
.c_out32(out_544),
.c_out33(out_545),
.c_out34(out_546),
.c_out35(out_547),
.c_out36(out_548),
.c_out37(out_549),
.c_out38(out_550),
.c_out39(out_551),
.c_out40(out_552),
.c_out41(out_553),
.c_out42(out_554),
.c_out43(out_555),
.c_out44(out_556),
.c_out45(out_557),
.c_out46(out_558),
.c_out47(out_559),
.c_out48(out_560),
.c_out49(out_561),
.c_out50(out_562),
.c_out51(out_563),
.c_out52(out_564),
.c_out53(out_565),
.c_out54(out_566),
.c_out55(out_567),
.c_out56(out_568),
.c_out57(out_569),
.c_out58(out_570),
.c_out59(out_571),
.c_out60(out_572),
.c_out61(out_573),
.c_out62(out_574),
.c_out63(out_575),
.c_out64(out_576),
.c_out65(out_577),
.c_out66(out_578),
.c_out67(out_579),
.c_out68(out_580),
.c_out69(out_581),
.c_out70(out_582),
.c_out71(out_583),
.c_out72(out_584),
.c_out73(out_585),
.c_out74(out_586),
.c_out75(out_587),
.c_out76(out_588),
.c_out77(out_589),
.c_out78(out_590),
.c_out79(out_591),
.c_out80(out_592),
.c_out81(out_593),
.c_out82(out_594),
.c_out83(out_595),
.c_out84(out_596),
.c_out85(out_597),
.c_out86(out_598),
.c_out87(out_599),
.c_out88(out_600),
.c_out89(out_601),
.c_out90(out_602),
.c_out91(out_603),
.c_out92(out_604),
.c_out93(out_605),
.c_out94(out_606),
.c_out95(out_607),
.c_out96(out_608),
.c_out97(out_609),
.c_out98(out_610),
.c_out99(out_611),
.c_out100(out_612),
.c_out101(out_613),
.c_out102(out_614),
.c_out103(out_615),
.c_out104(out_616),
.c_out105(out_617),
.c_out106(out_618),
.c_out107(out_619),
.c_out108(out_620),
.c_out109(out_621),
.c_out110(out_622),
.c_out111(out_623),
.c_out112(out_624),
.c_out113(out_625),
.c_out114(out_626),
.c_out115(out_627),
.c_out116(out_628),
.c_out117(out_629),
.c_out118(out_630),
.c_out119(out_631),
.c_out120(out_632),
.c_out121(out_633),
.c_out122(out_634),
.c_out123(out_635),
.c_out124(out_636),
.c_out125(out_637),
.c_out126(out_638),
.c_out127(out_639),
.c_out128(out_640),
.c_out129(out_641),
.c_out130(out_642),
.c_out131(out_643),
.c_out132(out_644),
.c_out133(out_645),
.c_out134(out_646),
.c_out135(out_647),
.c_out136(out_648),
.c_out137(out_649),
.c_out138(out_650),
.c_out139(out_651),
.c_out140(out_652),
.c_out141(out_653),
.c_out142(out_654),
.c_out143(out_655),
.c_out144(out_656),
.c_out145(out_657),
.c_out146(out_658),
.c_out147(out_659),
.c_out148(out_660),
.c_out149(out_661),
.c_out150(out_662),
.c_out151(out_663),
.c_out152(out_664),
.c_out153(out_665),
.c_out154(out_666),
.c_out155(out_667),
.c_out156(out_668),
.c_out157(out_669),
.c_out158(out_670),
.c_out159(out_671),
.c_out160(out_672),
.c_out161(out_673),
.c_out162(out_674),
.c_out163(out_675),
.c_out164(out_676),
.c_out165(out_677),
.c_out166(out_678),
.c_out167(out_679),
.c_out168(out_680),
.c_out169(out_681),
.c_out170(out_682),
.c_out171(out_683),
.c_out172(out_684),
.c_out173(out_685),
.c_out174(out_686),
.c_out175(out_687),
.c_out176(out_688),
.c_out177(out_689),
.c_out178(out_690),
.c_out179(out_691),
.c_out180(out_692),
.c_out181(out_693),
.c_out182(out_694),
.c_out183(out_695),
.c_out184(out_696),
.c_out185(out_697),
.c_out186(out_698),
.c_out187(out_699),
.c_out188(out_700),
.c_out189(out_701),
.c_out190(out_702),
.c_out191(out_703),
.c_out192(out_704),
.c_out193(out_705),
.c_out194(out_706),
.c_out195(out_707),
.c_out196(out_708),
.c_out197(out_709),
.c_out198(out_710),
.c_out199(out_711),
.c_out200(out_712),
.c_out201(out_713),
.c_out202(out_714),
.c_out203(out_715),
.c_out204(out_716),
.c_out205(out_717),
.c_out206(out_718),
.c_out207(out_719),
.c_out208(out_720),
.c_out209(out_721),
.c_out210(out_722),
.c_out211(out_723),
.c_out212(out_724),
.c_out213(out_725),
.c_out214(out_726),
.c_out215(out_727),
.c_out216(out_728),
.c_out217(out_729),
.c_out218(out_730),
.c_out219(out_731),
.c_out220(out_732),
.c_out221(out_733),
.c_out222(out_734),
.c_out223(out_735),
.c_out224(out_736),
.c_out225(out_737),
.c_out226(out_738),
.c_out227(out_739),
.c_out228(out_740),
.c_out229(out_741),
.c_out230(out_742),
.c_out231(out_743),
.c_out232(out_744),
.c_out233(out_745),
.c_out234(out_746),
.c_out235(out_747),
.c_out236(out_748),
.c_out237(out_749),
.c_out238(out_750),
.c_out239(out_751),
.c_out240(out_752),
.c_out241(out_753),
.c_out242(out_754),
.c_out243(out_755),
.c_out244(out_756),
.c_out245(out_757),
.c_out246(out_758),
.c_out247(out_759),
.c_out248(out_760),
.c_out249(out_761),
.c_out250(out_762),
.c_out251(out_763),
.c_out252(out_764),
.c_out253(out_765),
.c_out254(out_766),
.c_out255(out_767),
.c_out256(out_768),
.c_out257(out_769),
.c_out258(out_770),
.c_out259(out_771),
.c_out260(out_772),
.c_out261(out_773),
.c_out262(out_774),
.c_out263(out_775),
.c_out264(out_776),
.c_out265(out_777),
.c_out266(out_778),
.c_out267(out_779),
.c_out268(out_780),
.c_out269(out_781),
.c_out270(out_782),
.c_out271(out_783),
.c_out272(out_784),
.c_out273(out_785),
.c_out274(out_786),
.c_out275(out_787),
.c_out276(out_788),
.c_out277(out_789),
.c_out278(out_790),
.c_out279(out_791),
.c_out280(out_792),
.c_out281(out_793),
.c_out282(out_794),
.c_out283(out_795),
.c_out284(out_796),
.c_out285(out_797),
.c_out286(out_798),
.c_out287(out_799),
.c_out288(out_800),
.c_out289(out_801),
.c_out290(out_802),
.c_out291(out_803),
.c_out292(out_804),
.c_out293(out_805),
.c_out294(out_806),
.c_out295(out_807),
.c_out296(out_808),
.c_out297(out_809),
.c_out298(out_810),
.c_out299(out_811),
.c_out300(out_812),
.c_out301(out_813),
.c_out302(out_814),
.c_out303(out_815),
.c_out304(out_816),
.c_out305(out_817),
.c_out306(out_818),
.c_out307(out_819),
.c_out308(out_820),
.c_out309(out_821),
.c_out310(out_822),
.c_out311(out_823),
.c_out312(out_824),
.c_out313(out_825),
.c_out314(out_826),
.c_out315(out_827),
.c_out316(out_828),
.c_out317(out_829),
.c_out318(out_830),
.c_out319(out_831),
.c_out320(out_832),
.c_out321(out_833),
.c_out322(out_834),
.c_out323(out_835),
.c_out324(out_836),
.c_out325(out_837),
.c_out326(out_838),
.c_out327(out_839),
.c_out328(out_840),
.c_out329(out_841),
.c_out330(out_842),
.c_out331(out_843),
.c_out332(out_844),
.c_out333(out_845),
.c_out334(out_846),
.c_out335(out_847),
.c_out336(out_848),
.c_out337(out_849),
.c_out338(out_850),
.c_out339(out_851),
.c_out340(out_852),
.c_out341(out_853),
.c_out342(out_854),
.c_out343(out_855),
.c_out344(out_856),
.c_out345(out_857),
.c_out346(out_858),
.c_out347(out_859),
.c_out348(out_860),
.c_out349(out_861),
.c_out350(out_862),
.c_out351(out_863),
.c_out352(out_864),
.c_out353(out_865),
.c_out354(out_866),
.c_out355(out_867),
.c_out356(out_868),
.c_out357(out_869),
.c_out358(out_870),
.c_out359(out_871),
.c_out360(out_872),
.c_out361(out_873),
.c_out362(out_874),
.c_out363(out_875),
.c_out364(out_876),
.c_out365(out_877),
.c_out366(out_878),
.c_out367(out_879),
.c_out368(out_880),
.c_out369(out_881),
.c_out370(out_882),
.c_out371(out_883),
.c_out372(out_884),
.c_out373(out_885),
.c_out374(out_886),
.c_out375(out_887),
.c_out376(out_888),
.c_out377(out_889),
.c_out378(out_890),
.c_out379(out_891),
.c_out380(out_892),
.c_out381(out_893),
.c_out382(out_894),
.c_out383(out_895),
.c_out384(out_896),
.c_out385(out_897),
.c_out386(out_898),
.c_out387(out_899),
.c_out388(out_900),
.c_out389(out_901),
.c_out390(out_902),
.c_out391(out_903),
.c_out392(out_904),
.c_out393(out_905),
.c_out394(out_906),
.c_out395(out_907),
.c_out396(out_908),
.c_out397(out_909),
.c_out398(out_910),
.c_out399(out_911),
.c_out400(out_912),
.c_out401(out_913),
.c_out402(out_914),
.c_out403(out_915),
.c_out404(out_916),
.c_out405(out_917),
.c_out406(out_918),
.c_out407(out_919),
.c_out408(out_920),
.c_out409(out_921),
.c_out410(out_922),
.c_out411(out_923),
.c_out412(out_924),
.c_out413(out_925),
.c_out414(out_926),
.c_out415(out_927),
.c_out416(out_928),
.c_out417(out_929),
.c_out418(out_930),
.c_out419(out_931),
.c_out420(out_932),
.c_out421(out_933),
.c_out422(out_934),
.c_out423(out_935),
.c_out424(out_936),
.c_out425(out_937),
.c_out426(out_938),
.c_out427(out_939),
.c_out428(out_940),
.c_out429(out_941),
.c_out430(out_942),
.c_out431(out_943),
.c_out432(out_944),
.c_out433(out_945),
.c_out434(out_946),
.c_out435(out_947),
.c_out436(out_948),
.c_out437(out_949),
.c_out438(out_950),
.c_out439(out_951),
.c_out440(out_952),
.c_out441(out_953),
.c_out442(out_954),
.c_out443(out_955),
.c_out444(out_956),
.c_out445(out_957),
.c_out446(out_958),
.c_out447(out_959),
.c_out448(out_960),
.c_out449(out_961),
.c_out450(out_962),
.c_out451(out_963),
.c_out452(out_964),
.c_out453(out_965),
.c_out454(out_966),
.c_out455(out_967),
.c_out456(out_968),
.c_out457(out_969),
.c_out458(out_970),
.c_out459(out_971),
.c_out460(out_972),
.c_out461(out_973),
.c_out462(out_974),
.c_out463(out_975),
.c_out464(out_976),
.c_out465(out_977),
.c_out466(out_978),
.c_out467(out_979),
.c_out468(out_980),
.c_out469(out_981),
.c_out470(out_982),
.c_out471(out_983),
.c_out472(out_984),
.c_out473(out_985),
.c_out474(out_986),
.c_out475(out_987),
.c_out476(out_988),
.c_out477(out_989),
.c_out478(out_990),
.c_out479(out_991),
.c_out480(out_992),
.c_out481(out_993),
.c_out482(out_994),
.c_out483(out_995),
.c_out484(out_996),
.c_out485(out_997),
.c_out486(out_998),
.c_out487(out_999),
.c_out488(out_1000),
.c_out489(out_1001),
.c_out490(out_1002),
.c_out491(out_1003),
.c_out492(out_1004),
.c_out493(out_1005),
.c_out494(out_1006),
.c_out495(out_1007),
.c_out496(out_1008),
.c_out497(out_1009),
.c_out498(out_1010),
.c_out499(out_1011),
.c_out500(out_1012),
.c_out501(out_1013),
.c_out502(out_1014),
.c_out503(out_1015),
.c_out504(out_1016),
.c_out505(out_1017),
.c_out506(out_1018),
.c_out507(out_1019),
.c_out508(out_1020),
.c_out509(out_1021),
.c_out510(out_1022),
.c_out511(out_1023));
SA128 SA128_2 (.clk(clk),.rstn(rstn),.activation(act_1),.weight(weight0_2),.out_act(act2_3),.out_weight(outweight_0),.control(control),.c_out0(out_1024),
.c_out1(out_1025),
.c_out2(out_1026),
.c_out3(out_1027),
.c_out4(out_1028),
.c_out5(out_1029),
.c_out6(out_1030),
.c_out7(out_1031),
.c_out8(out_1032),
.c_out9(out_1033),
.c_out10(out_1034),
.c_out11(out_1035),
.c_out12(out_1036),
.c_out13(out_1037),
.c_out14(out_1038),
.c_out15(out_1039),
.c_out16(out_1040),
.c_out17(out_1041),
.c_out18(out_1042),
.c_out19(out_1043),
.c_out20(out_1044),
.c_out21(out_1045),
.c_out22(out_1046),
.c_out23(out_1047),
.c_out24(out_1048),
.c_out25(out_1049),
.c_out26(out_1050),
.c_out27(out_1051),
.c_out28(out_1052),
.c_out29(out_1053),
.c_out30(out_1054),
.c_out31(out_1055),
.c_out32(out_1056),
.c_out33(out_1057),
.c_out34(out_1058),
.c_out35(out_1059),
.c_out36(out_1060),
.c_out37(out_1061),
.c_out38(out_1062),
.c_out39(out_1063),
.c_out40(out_1064),
.c_out41(out_1065),
.c_out42(out_1066),
.c_out43(out_1067),
.c_out44(out_1068),
.c_out45(out_1069),
.c_out46(out_1070),
.c_out47(out_1071),
.c_out48(out_1072),
.c_out49(out_1073),
.c_out50(out_1074),
.c_out51(out_1075),
.c_out52(out_1076),
.c_out53(out_1077),
.c_out54(out_1078),
.c_out55(out_1079),
.c_out56(out_1080),
.c_out57(out_1081),
.c_out58(out_1082),
.c_out59(out_1083),
.c_out60(out_1084),
.c_out61(out_1085),
.c_out62(out_1086),
.c_out63(out_1087),
.c_out64(out_1088),
.c_out65(out_1089),
.c_out66(out_1090),
.c_out67(out_1091),
.c_out68(out_1092),
.c_out69(out_1093),
.c_out70(out_1094),
.c_out71(out_1095),
.c_out72(out_1096),
.c_out73(out_1097),
.c_out74(out_1098),
.c_out75(out_1099),
.c_out76(out_1100),
.c_out77(out_1101),
.c_out78(out_1102),
.c_out79(out_1103),
.c_out80(out_1104),
.c_out81(out_1105),
.c_out82(out_1106),
.c_out83(out_1107),
.c_out84(out_1108),
.c_out85(out_1109),
.c_out86(out_1110),
.c_out87(out_1111),
.c_out88(out_1112),
.c_out89(out_1113),
.c_out90(out_1114),
.c_out91(out_1115),
.c_out92(out_1116),
.c_out93(out_1117),
.c_out94(out_1118),
.c_out95(out_1119),
.c_out96(out_1120),
.c_out97(out_1121),
.c_out98(out_1122),
.c_out99(out_1123),
.c_out100(out_1124),
.c_out101(out_1125),
.c_out102(out_1126),
.c_out103(out_1127),
.c_out104(out_1128),
.c_out105(out_1129),
.c_out106(out_1130),
.c_out107(out_1131),
.c_out108(out_1132),
.c_out109(out_1133),
.c_out110(out_1134),
.c_out111(out_1135),
.c_out112(out_1136),
.c_out113(out_1137),
.c_out114(out_1138),
.c_out115(out_1139),
.c_out116(out_1140),
.c_out117(out_1141),
.c_out118(out_1142),
.c_out119(out_1143),
.c_out120(out_1144),
.c_out121(out_1145),
.c_out122(out_1146),
.c_out123(out_1147),
.c_out124(out_1148),
.c_out125(out_1149),
.c_out126(out_1150),
.c_out127(out_1151),
.c_out128(out_1152),
.c_out129(out_1153),
.c_out130(out_1154),
.c_out131(out_1155),
.c_out132(out_1156),
.c_out133(out_1157),
.c_out134(out_1158),
.c_out135(out_1159),
.c_out136(out_1160),
.c_out137(out_1161),
.c_out138(out_1162),
.c_out139(out_1163),
.c_out140(out_1164),
.c_out141(out_1165),
.c_out142(out_1166),
.c_out143(out_1167),
.c_out144(out_1168),
.c_out145(out_1169),
.c_out146(out_1170),
.c_out147(out_1171),
.c_out148(out_1172),
.c_out149(out_1173),
.c_out150(out_1174),
.c_out151(out_1175),
.c_out152(out_1176),
.c_out153(out_1177),
.c_out154(out_1178),
.c_out155(out_1179),
.c_out156(out_1180),
.c_out157(out_1181),
.c_out158(out_1182),
.c_out159(out_1183),
.c_out160(out_1184),
.c_out161(out_1185),
.c_out162(out_1186),
.c_out163(out_1187),
.c_out164(out_1188),
.c_out165(out_1189),
.c_out166(out_1190),
.c_out167(out_1191),
.c_out168(out_1192),
.c_out169(out_1193),
.c_out170(out_1194),
.c_out171(out_1195),
.c_out172(out_1196),
.c_out173(out_1197),
.c_out174(out_1198),
.c_out175(out_1199),
.c_out176(out_1200),
.c_out177(out_1201),
.c_out178(out_1202),
.c_out179(out_1203),
.c_out180(out_1204),
.c_out181(out_1205),
.c_out182(out_1206),
.c_out183(out_1207),
.c_out184(out_1208),
.c_out185(out_1209),
.c_out186(out_1210),
.c_out187(out_1211),
.c_out188(out_1212),
.c_out189(out_1213),
.c_out190(out_1214),
.c_out191(out_1215),
.c_out192(out_1216),
.c_out193(out_1217),
.c_out194(out_1218),
.c_out195(out_1219),
.c_out196(out_1220),
.c_out197(out_1221),
.c_out198(out_1222),
.c_out199(out_1223),
.c_out200(out_1224),
.c_out201(out_1225),
.c_out202(out_1226),
.c_out203(out_1227),
.c_out204(out_1228),
.c_out205(out_1229),
.c_out206(out_1230),
.c_out207(out_1231),
.c_out208(out_1232),
.c_out209(out_1233),
.c_out210(out_1234),
.c_out211(out_1235),
.c_out212(out_1236),
.c_out213(out_1237),
.c_out214(out_1238),
.c_out215(out_1239),
.c_out216(out_1240),
.c_out217(out_1241),
.c_out218(out_1242),
.c_out219(out_1243),
.c_out220(out_1244),
.c_out221(out_1245),
.c_out222(out_1246),
.c_out223(out_1247),
.c_out224(out_1248),
.c_out225(out_1249),
.c_out226(out_1250),
.c_out227(out_1251),
.c_out228(out_1252),
.c_out229(out_1253),
.c_out230(out_1254),
.c_out231(out_1255),
.c_out232(out_1256),
.c_out233(out_1257),
.c_out234(out_1258),
.c_out235(out_1259),
.c_out236(out_1260),
.c_out237(out_1261),
.c_out238(out_1262),
.c_out239(out_1263),
.c_out240(out_1264),
.c_out241(out_1265),
.c_out242(out_1266),
.c_out243(out_1267),
.c_out244(out_1268),
.c_out245(out_1269),
.c_out246(out_1270),
.c_out247(out_1271),
.c_out248(out_1272),
.c_out249(out_1273),
.c_out250(out_1274),
.c_out251(out_1275),
.c_out252(out_1276),
.c_out253(out_1277),
.c_out254(out_1278),
.c_out255(out_1279),
.c_out256(out_1280),
.c_out257(out_1281),
.c_out258(out_1282),
.c_out259(out_1283),
.c_out260(out_1284),
.c_out261(out_1285),
.c_out262(out_1286),
.c_out263(out_1287),
.c_out264(out_1288),
.c_out265(out_1289),
.c_out266(out_1290),
.c_out267(out_1291),
.c_out268(out_1292),
.c_out269(out_1293),
.c_out270(out_1294),
.c_out271(out_1295),
.c_out272(out_1296),
.c_out273(out_1297),
.c_out274(out_1298),
.c_out275(out_1299),
.c_out276(out_1300),
.c_out277(out_1301),
.c_out278(out_1302),
.c_out279(out_1303),
.c_out280(out_1304),
.c_out281(out_1305),
.c_out282(out_1306),
.c_out283(out_1307),
.c_out284(out_1308),
.c_out285(out_1309),
.c_out286(out_1310),
.c_out287(out_1311),
.c_out288(out_1312),
.c_out289(out_1313),
.c_out290(out_1314),
.c_out291(out_1315),
.c_out292(out_1316),
.c_out293(out_1317),
.c_out294(out_1318),
.c_out295(out_1319),
.c_out296(out_1320),
.c_out297(out_1321),
.c_out298(out_1322),
.c_out299(out_1323),
.c_out300(out_1324),
.c_out301(out_1325),
.c_out302(out_1326),
.c_out303(out_1327),
.c_out304(out_1328),
.c_out305(out_1329),
.c_out306(out_1330),
.c_out307(out_1331),
.c_out308(out_1332),
.c_out309(out_1333),
.c_out310(out_1334),
.c_out311(out_1335),
.c_out312(out_1336),
.c_out313(out_1337),
.c_out314(out_1338),
.c_out315(out_1339),
.c_out316(out_1340),
.c_out317(out_1341),
.c_out318(out_1342),
.c_out319(out_1343),
.c_out320(out_1344),
.c_out321(out_1345),
.c_out322(out_1346),
.c_out323(out_1347),
.c_out324(out_1348),
.c_out325(out_1349),
.c_out326(out_1350),
.c_out327(out_1351),
.c_out328(out_1352),
.c_out329(out_1353),
.c_out330(out_1354),
.c_out331(out_1355),
.c_out332(out_1356),
.c_out333(out_1357),
.c_out334(out_1358),
.c_out335(out_1359),
.c_out336(out_1360),
.c_out337(out_1361),
.c_out338(out_1362),
.c_out339(out_1363),
.c_out340(out_1364),
.c_out341(out_1365),
.c_out342(out_1366),
.c_out343(out_1367),
.c_out344(out_1368),
.c_out345(out_1369),
.c_out346(out_1370),
.c_out347(out_1371),
.c_out348(out_1372),
.c_out349(out_1373),
.c_out350(out_1374),
.c_out351(out_1375),
.c_out352(out_1376),
.c_out353(out_1377),
.c_out354(out_1378),
.c_out355(out_1379),
.c_out356(out_1380),
.c_out357(out_1381),
.c_out358(out_1382),
.c_out359(out_1383),
.c_out360(out_1384),
.c_out361(out_1385),
.c_out362(out_1386),
.c_out363(out_1387),
.c_out364(out_1388),
.c_out365(out_1389),
.c_out366(out_1390),
.c_out367(out_1391),
.c_out368(out_1392),
.c_out369(out_1393),
.c_out370(out_1394),
.c_out371(out_1395),
.c_out372(out_1396),
.c_out373(out_1397),
.c_out374(out_1398),
.c_out375(out_1399),
.c_out376(out_1400),
.c_out377(out_1401),
.c_out378(out_1402),
.c_out379(out_1403),
.c_out380(out_1404),
.c_out381(out_1405),
.c_out382(out_1406),
.c_out383(out_1407),
.c_out384(out_1408),
.c_out385(out_1409),
.c_out386(out_1410),
.c_out387(out_1411),
.c_out388(out_1412),
.c_out389(out_1413),
.c_out390(out_1414),
.c_out391(out_1415),
.c_out392(out_1416),
.c_out393(out_1417),
.c_out394(out_1418),
.c_out395(out_1419),
.c_out396(out_1420),
.c_out397(out_1421),
.c_out398(out_1422),
.c_out399(out_1423),
.c_out400(out_1424),
.c_out401(out_1425),
.c_out402(out_1426),
.c_out403(out_1427),
.c_out404(out_1428),
.c_out405(out_1429),
.c_out406(out_1430),
.c_out407(out_1431),
.c_out408(out_1432),
.c_out409(out_1433),
.c_out410(out_1434),
.c_out411(out_1435),
.c_out412(out_1436),
.c_out413(out_1437),
.c_out414(out_1438),
.c_out415(out_1439),
.c_out416(out_1440),
.c_out417(out_1441),
.c_out418(out_1442),
.c_out419(out_1443),
.c_out420(out_1444),
.c_out421(out_1445),
.c_out422(out_1446),
.c_out423(out_1447),
.c_out424(out_1448),
.c_out425(out_1449),
.c_out426(out_1450),
.c_out427(out_1451),
.c_out428(out_1452),
.c_out429(out_1453),
.c_out430(out_1454),
.c_out431(out_1455),
.c_out432(out_1456),
.c_out433(out_1457),
.c_out434(out_1458),
.c_out435(out_1459),
.c_out436(out_1460),
.c_out437(out_1461),
.c_out438(out_1462),
.c_out439(out_1463),
.c_out440(out_1464),
.c_out441(out_1465),
.c_out442(out_1466),
.c_out443(out_1467),
.c_out444(out_1468),
.c_out445(out_1469),
.c_out446(out_1470),
.c_out447(out_1471),
.c_out448(out_1472),
.c_out449(out_1473),
.c_out450(out_1474),
.c_out451(out_1475),
.c_out452(out_1476),
.c_out453(out_1477),
.c_out454(out_1478),
.c_out455(out_1479),
.c_out456(out_1480),
.c_out457(out_1481),
.c_out458(out_1482),
.c_out459(out_1483),
.c_out460(out_1484),
.c_out461(out_1485),
.c_out462(out_1486),
.c_out463(out_1487),
.c_out464(out_1488),
.c_out465(out_1489),
.c_out466(out_1490),
.c_out467(out_1491),
.c_out468(out_1492),
.c_out469(out_1493),
.c_out470(out_1494),
.c_out471(out_1495),
.c_out472(out_1496),
.c_out473(out_1497),
.c_out474(out_1498),
.c_out475(out_1499),
.c_out476(out_1500),
.c_out477(out_1501),
.c_out478(out_1502),
.c_out479(out_1503),
.c_out480(out_1504),
.c_out481(out_1505),
.c_out482(out_1506),
.c_out483(out_1507),
.c_out484(out_1508),
.c_out485(out_1509),
.c_out486(out_1510),
.c_out487(out_1511),
.c_out488(out_1512),
.c_out489(out_1513),
.c_out490(out_1514),
.c_out491(out_1515),
.c_out492(out_1516),
.c_out493(out_1517),
.c_out494(out_1518),
.c_out495(out_1519),
.c_out496(out_1520),
.c_out497(out_1521),
.c_out498(out_1522),
.c_out499(out_1523),
.c_out500(out_1524),
.c_out501(out_1525),
.c_out502(out_1526),
.c_out503(out_1527),
.c_out504(out_1528),
.c_out505(out_1529),
.c_out506(out_1530),
.c_out507(out_1531),
.c_out508(out_1532),
.c_out509(out_1533),
.c_out510(out_1534),
.c_out511(out_1535));
SA128 SA128_3 (.clk(clk),.rstn(rstn),.activation(act2_3),.weight(weight1_3),.out_act(outact_1),.out_weight(outweight_1),.control(control),.c_out0(out_1536),
.c_out1(out_1537),
.c_out2(out_1538),
.c_out3(out_1539),
.c_out4(out_1540),
.c_out5(out_1541),
.c_out6(out_1542),
.c_out7(out_1543),
.c_out8(out_1544),
.c_out9(out_1545),
.c_out10(out_1546),
.c_out11(out_1547),
.c_out12(out_1548),
.c_out13(out_1549),
.c_out14(out_1550),
.c_out15(out_1551),
.c_out16(out_1552),
.c_out17(out_1553),
.c_out18(out_1554),
.c_out19(out_1555),
.c_out20(out_1556),
.c_out21(out_1557),
.c_out22(out_1558),
.c_out23(out_1559),
.c_out24(out_1560),
.c_out25(out_1561),
.c_out26(out_1562),
.c_out27(out_1563),
.c_out28(out_1564),
.c_out29(out_1565),
.c_out30(out_1566),
.c_out31(out_1567),
.c_out32(out_1568),
.c_out33(out_1569),
.c_out34(out_1570),
.c_out35(out_1571),
.c_out36(out_1572),
.c_out37(out_1573),
.c_out38(out_1574),
.c_out39(out_1575),
.c_out40(out_1576),
.c_out41(out_1577),
.c_out42(out_1578),
.c_out43(out_1579),
.c_out44(out_1580),
.c_out45(out_1581),
.c_out46(out_1582),
.c_out47(out_1583),
.c_out48(out_1584),
.c_out49(out_1585),
.c_out50(out_1586),
.c_out51(out_1587),
.c_out52(out_1588),
.c_out53(out_1589),
.c_out54(out_1590),
.c_out55(out_1591),
.c_out56(out_1592),
.c_out57(out_1593),
.c_out58(out_1594),
.c_out59(out_1595),
.c_out60(out_1596),
.c_out61(out_1597),
.c_out62(out_1598),
.c_out63(out_1599),
.c_out64(out_1600),
.c_out65(out_1601),
.c_out66(out_1602),
.c_out67(out_1603),
.c_out68(out_1604),
.c_out69(out_1605),
.c_out70(out_1606),
.c_out71(out_1607),
.c_out72(out_1608),
.c_out73(out_1609),
.c_out74(out_1610),
.c_out75(out_1611),
.c_out76(out_1612),
.c_out77(out_1613),
.c_out78(out_1614),
.c_out79(out_1615),
.c_out80(out_1616),
.c_out81(out_1617),
.c_out82(out_1618),
.c_out83(out_1619),
.c_out84(out_1620),
.c_out85(out_1621),
.c_out86(out_1622),
.c_out87(out_1623),
.c_out88(out_1624),
.c_out89(out_1625),
.c_out90(out_1626),
.c_out91(out_1627),
.c_out92(out_1628),
.c_out93(out_1629),
.c_out94(out_1630),
.c_out95(out_1631),
.c_out96(out_1632),
.c_out97(out_1633),
.c_out98(out_1634),
.c_out99(out_1635),
.c_out100(out_1636),
.c_out101(out_1637),
.c_out102(out_1638),
.c_out103(out_1639),
.c_out104(out_1640),
.c_out105(out_1641),
.c_out106(out_1642),
.c_out107(out_1643),
.c_out108(out_1644),
.c_out109(out_1645),
.c_out110(out_1646),
.c_out111(out_1647),
.c_out112(out_1648),
.c_out113(out_1649),
.c_out114(out_1650),
.c_out115(out_1651),
.c_out116(out_1652),
.c_out117(out_1653),
.c_out118(out_1654),
.c_out119(out_1655),
.c_out120(out_1656),
.c_out121(out_1657),
.c_out122(out_1658),
.c_out123(out_1659),
.c_out124(out_1660),
.c_out125(out_1661),
.c_out126(out_1662),
.c_out127(out_1663),
.c_out128(out_1664),
.c_out129(out_1665),
.c_out130(out_1666),
.c_out131(out_1667),
.c_out132(out_1668),
.c_out133(out_1669),
.c_out134(out_1670),
.c_out135(out_1671),
.c_out136(out_1672),
.c_out137(out_1673),
.c_out138(out_1674),
.c_out139(out_1675),
.c_out140(out_1676),
.c_out141(out_1677),
.c_out142(out_1678),
.c_out143(out_1679),
.c_out144(out_1680),
.c_out145(out_1681),
.c_out146(out_1682),
.c_out147(out_1683),
.c_out148(out_1684),
.c_out149(out_1685),
.c_out150(out_1686),
.c_out151(out_1687),
.c_out152(out_1688),
.c_out153(out_1689),
.c_out154(out_1690),
.c_out155(out_1691),
.c_out156(out_1692),
.c_out157(out_1693),
.c_out158(out_1694),
.c_out159(out_1695),
.c_out160(out_1696),
.c_out161(out_1697),
.c_out162(out_1698),
.c_out163(out_1699),
.c_out164(out_1700),
.c_out165(out_1701),
.c_out166(out_1702),
.c_out167(out_1703),
.c_out168(out_1704),
.c_out169(out_1705),
.c_out170(out_1706),
.c_out171(out_1707),
.c_out172(out_1708),
.c_out173(out_1709),
.c_out174(out_1710),
.c_out175(out_1711),
.c_out176(out_1712),
.c_out177(out_1713),
.c_out178(out_1714),
.c_out179(out_1715),
.c_out180(out_1716),
.c_out181(out_1717),
.c_out182(out_1718),
.c_out183(out_1719),
.c_out184(out_1720),
.c_out185(out_1721),
.c_out186(out_1722),
.c_out187(out_1723),
.c_out188(out_1724),
.c_out189(out_1725),
.c_out190(out_1726),
.c_out191(out_1727),
.c_out192(out_1728),
.c_out193(out_1729),
.c_out194(out_1730),
.c_out195(out_1731),
.c_out196(out_1732),
.c_out197(out_1733),
.c_out198(out_1734),
.c_out199(out_1735),
.c_out200(out_1736),
.c_out201(out_1737),
.c_out202(out_1738),
.c_out203(out_1739),
.c_out204(out_1740),
.c_out205(out_1741),
.c_out206(out_1742),
.c_out207(out_1743),
.c_out208(out_1744),
.c_out209(out_1745),
.c_out210(out_1746),
.c_out211(out_1747),
.c_out212(out_1748),
.c_out213(out_1749),
.c_out214(out_1750),
.c_out215(out_1751),
.c_out216(out_1752),
.c_out217(out_1753),
.c_out218(out_1754),
.c_out219(out_1755),
.c_out220(out_1756),
.c_out221(out_1757),
.c_out222(out_1758),
.c_out223(out_1759),
.c_out224(out_1760),
.c_out225(out_1761),
.c_out226(out_1762),
.c_out227(out_1763),
.c_out228(out_1764),
.c_out229(out_1765),
.c_out230(out_1766),
.c_out231(out_1767),
.c_out232(out_1768),
.c_out233(out_1769),
.c_out234(out_1770),
.c_out235(out_1771),
.c_out236(out_1772),
.c_out237(out_1773),
.c_out238(out_1774),
.c_out239(out_1775),
.c_out240(out_1776),
.c_out241(out_1777),
.c_out242(out_1778),
.c_out243(out_1779),
.c_out244(out_1780),
.c_out245(out_1781),
.c_out246(out_1782),
.c_out247(out_1783),
.c_out248(out_1784),
.c_out249(out_1785),
.c_out250(out_1786),
.c_out251(out_1787),
.c_out252(out_1788),
.c_out253(out_1789),
.c_out254(out_1790),
.c_out255(out_1791),
.c_out256(out_1792),
.c_out257(out_1793),
.c_out258(out_1794),
.c_out259(out_1795),
.c_out260(out_1796),
.c_out261(out_1797),
.c_out262(out_1798),
.c_out263(out_1799),
.c_out264(out_1800),
.c_out265(out_1801),
.c_out266(out_1802),
.c_out267(out_1803),
.c_out268(out_1804),
.c_out269(out_1805),
.c_out270(out_1806),
.c_out271(out_1807),
.c_out272(out_1808),
.c_out273(out_1809),
.c_out274(out_1810),
.c_out275(out_1811),
.c_out276(out_1812),
.c_out277(out_1813),
.c_out278(out_1814),
.c_out279(out_1815),
.c_out280(out_1816),
.c_out281(out_1817),
.c_out282(out_1818),
.c_out283(out_1819),
.c_out284(out_1820),
.c_out285(out_1821),
.c_out286(out_1822),
.c_out287(out_1823),
.c_out288(out_1824),
.c_out289(out_1825),
.c_out290(out_1826),
.c_out291(out_1827),
.c_out292(out_1828),
.c_out293(out_1829),
.c_out294(out_1830),
.c_out295(out_1831),
.c_out296(out_1832),
.c_out297(out_1833),
.c_out298(out_1834),
.c_out299(out_1835),
.c_out300(out_1836),
.c_out301(out_1837),
.c_out302(out_1838),
.c_out303(out_1839),
.c_out304(out_1840),
.c_out305(out_1841),
.c_out306(out_1842),
.c_out307(out_1843),
.c_out308(out_1844),
.c_out309(out_1845),
.c_out310(out_1846),
.c_out311(out_1847),
.c_out312(out_1848),
.c_out313(out_1849),
.c_out314(out_1850),
.c_out315(out_1851),
.c_out316(out_1852),
.c_out317(out_1853),
.c_out318(out_1854),
.c_out319(out_1855),
.c_out320(out_1856),
.c_out321(out_1857),
.c_out322(out_1858),
.c_out323(out_1859),
.c_out324(out_1860),
.c_out325(out_1861),
.c_out326(out_1862),
.c_out327(out_1863),
.c_out328(out_1864),
.c_out329(out_1865),
.c_out330(out_1866),
.c_out331(out_1867),
.c_out332(out_1868),
.c_out333(out_1869),
.c_out334(out_1870),
.c_out335(out_1871),
.c_out336(out_1872),
.c_out337(out_1873),
.c_out338(out_1874),
.c_out339(out_1875),
.c_out340(out_1876),
.c_out341(out_1877),
.c_out342(out_1878),
.c_out343(out_1879),
.c_out344(out_1880),
.c_out345(out_1881),
.c_out346(out_1882),
.c_out347(out_1883),
.c_out348(out_1884),
.c_out349(out_1885),
.c_out350(out_1886),
.c_out351(out_1887),
.c_out352(out_1888),
.c_out353(out_1889),
.c_out354(out_1890),
.c_out355(out_1891),
.c_out356(out_1892),
.c_out357(out_1893),
.c_out358(out_1894),
.c_out359(out_1895),
.c_out360(out_1896),
.c_out361(out_1897),
.c_out362(out_1898),
.c_out363(out_1899),
.c_out364(out_1900),
.c_out365(out_1901),
.c_out366(out_1902),
.c_out367(out_1903),
.c_out368(out_1904),
.c_out369(out_1905),
.c_out370(out_1906),
.c_out371(out_1907),
.c_out372(out_1908),
.c_out373(out_1909),
.c_out374(out_1910),
.c_out375(out_1911),
.c_out376(out_1912),
.c_out377(out_1913),
.c_out378(out_1914),
.c_out379(out_1915),
.c_out380(out_1916),
.c_out381(out_1917),
.c_out382(out_1918),
.c_out383(out_1919),
.c_out384(out_1920),
.c_out385(out_1921),
.c_out386(out_1922),
.c_out387(out_1923),
.c_out388(out_1924),
.c_out389(out_1925),
.c_out390(out_1926),
.c_out391(out_1927),
.c_out392(out_1928),
.c_out393(out_1929),
.c_out394(out_1930),
.c_out395(out_1931),
.c_out396(out_1932),
.c_out397(out_1933),
.c_out398(out_1934),
.c_out399(out_1935),
.c_out400(out_1936),
.c_out401(out_1937),
.c_out402(out_1938),
.c_out403(out_1939),
.c_out404(out_1940),
.c_out405(out_1941),
.c_out406(out_1942),
.c_out407(out_1943),
.c_out408(out_1944),
.c_out409(out_1945),
.c_out410(out_1946),
.c_out411(out_1947),
.c_out412(out_1948),
.c_out413(out_1949),
.c_out414(out_1950),
.c_out415(out_1951),
.c_out416(out_1952),
.c_out417(out_1953),
.c_out418(out_1954),
.c_out419(out_1955),
.c_out420(out_1956),
.c_out421(out_1957),
.c_out422(out_1958),
.c_out423(out_1959),
.c_out424(out_1960),
.c_out425(out_1961),
.c_out426(out_1962),
.c_out427(out_1963),
.c_out428(out_1964),
.c_out429(out_1965),
.c_out430(out_1966),
.c_out431(out_1967),
.c_out432(out_1968),
.c_out433(out_1969),
.c_out434(out_1970),
.c_out435(out_1971),
.c_out436(out_1972),
.c_out437(out_1973),
.c_out438(out_1974),
.c_out439(out_1975),
.c_out440(out_1976),
.c_out441(out_1977),
.c_out442(out_1978),
.c_out443(out_1979),
.c_out444(out_1980),
.c_out445(out_1981),
.c_out446(out_1982),
.c_out447(out_1983),
.c_out448(out_1984),
.c_out449(out_1985),
.c_out450(out_1986),
.c_out451(out_1987),
.c_out452(out_1988),
.c_out453(out_1989),
.c_out454(out_1990),
.c_out455(out_1991),
.c_out456(out_1992),
.c_out457(out_1993),
.c_out458(out_1994),
.c_out459(out_1995),
.c_out460(out_1996),
.c_out461(out_1997),
.c_out462(out_1998),
.c_out463(out_1999),
.c_out464(out_2000),
.c_out465(out_2001),
.c_out466(out_2002),
.c_out467(out_2003),
.c_out468(out_2004),
.c_out469(out_2005),
.c_out470(out_2006),
.c_out471(out_2007),
.c_out472(out_2008),
.c_out473(out_2009),
.c_out474(out_2010),
.c_out475(out_2011),
.c_out476(out_2012),
.c_out477(out_2013),
.c_out478(out_2014),
.c_out479(out_2015),
.c_out480(out_2016),
.c_out481(out_2017),
.c_out482(out_2018),
.c_out483(out_2019),
.c_out484(out_2020),
.c_out485(out_2021),
.c_out486(out_2022),
.c_out487(out_2023),
.c_out488(out_2024),
.c_out489(out_2025),
.c_out490(out_2026),
.c_out491(out_2027),
.c_out492(out_2028),
.c_out493(out_2029),
.c_out494(out_2030),
.c_out495(out_2031),
.c_out496(out_2032),
.c_out497(out_2033),
.c_out498(out_2034),
.c_out499(out_2035),
.c_out500(out_2036),
.c_out501(out_2037),
.c_out502(out_2038),
.c_out503(out_2039),
.c_out504(out_2040),
.c_out505(out_2041),
.c_out506(out_2042),
.c_out507(out_2043),
.c_out508(out_2044),
.c_out509(out_2045),
.c_out510(out_2046),
.c_out511(out_2047));

assign out_act = {outact_0,outact_1};
assign out_weight = {outweight_0,outweight_1};

assign c_out0 = out_0;
assign c_out1 = out_1;
assign c_out2 = out_2;
assign c_out3 = out_3;
assign c_out4 = out_4;
assign c_out5 = out_5;
assign c_out6 = out_6;
assign c_out7 = out_7;
assign c_out8 = out_8;
assign c_out9 = out_9;
assign c_out10 = out_10;
assign c_out11 = out_11;
assign c_out12 = out_12;
assign c_out13 = out_13;
assign c_out14 = out_14;
assign c_out15 = out_15;
assign c_out16 = out_16;
assign c_out17 = out_17;
assign c_out18 = out_18;
assign c_out19 = out_19;
assign c_out20 = out_20;
assign c_out21 = out_21;
assign c_out22 = out_22;
assign c_out23 = out_23;
assign c_out24 = out_24;
assign c_out25 = out_25;
assign c_out26 = out_26;
assign c_out27 = out_27;
assign c_out28 = out_28;
assign c_out29 = out_29;
assign c_out30 = out_30;
assign c_out31 = out_31;
assign c_out32 = out_32;
assign c_out33 = out_33;
assign c_out34 = out_34;
assign c_out35 = out_35;
assign c_out36 = out_36;
assign c_out37 = out_37;
assign c_out38 = out_38;
assign c_out39 = out_39;
assign c_out40 = out_40;
assign c_out41 = out_41;
assign c_out42 = out_42;
assign c_out43 = out_43;
assign c_out44 = out_44;
assign c_out45 = out_45;
assign c_out46 = out_46;
assign c_out47 = out_47;
assign c_out48 = out_48;
assign c_out49 = out_49;
assign c_out50 = out_50;
assign c_out51 = out_51;
assign c_out52 = out_52;
assign c_out53 = out_53;
assign c_out54 = out_54;
assign c_out55 = out_55;
assign c_out56 = out_56;
assign c_out57 = out_57;
assign c_out58 = out_58;
assign c_out59 = out_59;
assign c_out60 = out_60;
assign c_out61 = out_61;
assign c_out62 = out_62;
assign c_out63 = out_63;
assign c_out64 = out_64;
assign c_out65 = out_65;
assign c_out66 = out_66;
assign c_out67 = out_67;
assign c_out68 = out_68;
assign c_out69 = out_69;
assign c_out70 = out_70;
assign c_out71 = out_71;
assign c_out72 = out_72;
assign c_out73 = out_73;
assign c_out74 = out_74;
assign c_out75 = out_75;
assign c_out76 = out_76;
assign c_out77 = out_77;
assign c_out78 = out_78;
assign c_out79 = out_79;
assign c_out80 = out_80;
assign c_out81 = out_81;
assign c_out82 = out_82;
assign c_out83 = out_83;
assign c_out84 = out_84;
assign c_out85 = out_85;
assign c_out86 = out_86;
assign c_out87 = out_87;
assign c_out88 = out_88;
assign c_out89 = out_89;
assign c_out90 = out_90;
assign c_out91 = out_91;
assign c_out92 = out_92;
assign c_out93 = out_93;
assign c_out94 = out_94;
assign c_out95 = out_95;
assign c_out96 = out_96;
assign c_out97 = out_97;
assign c_out98 = out_98;
assign c_out99 = out_99;
assign c_out100 = out_100;
assign c_out101 = out_101;
assign c_out102 = out_102;
assign c_out103 = out_103;
assign c_out104 = out_104;
assign c_out105 = out_105;
assign c_out106 = out_106;
assign c_out107 = out_107;
assign c_out108 = out_108;
assign c_out109 = out_109;
assign c_out110 = out_110;
assign c_out111 = out_111;
assign c_out112 = out_112;
assign c_out113 = out_113;
assign c_out114 = out_114;
assign c_out115 = out_115;
assign c_out116 = out_116;
assign c_out117 = out_117;
assign c_out118 = out_118;
assign c_out119 = out_119;
assign c_out120 = out_120;
assign c_out121 = out_121;
assign c_out122 = out_122;
assign c_out123 = out_123;
assign c_out124 = out_124;
assign c_out125 = out_125;
assign c_out126 = out_126;
assign c_out127 = out_127;
assign c_out128 = out_128;
assign c_out129 = out_129;
assign c_out130 = out_130;
assign c_out131 = out_131;
assign c_out132 = out_132;
assign c_out133 = out_133;
assign c_out134 = out_134;
assign c_out135 = out_135;
assign c_out136 = out_136;
assign c_out137 = out_137;
assign c_out138 = out_138;
assign c_out139 = out_139;
assign c_out140 = out_140;
assign c_out141 = out_141;
assign c_out142 = out_142;
assign c_out143 = out_143;
assign c_out144 = out_144;
assign c_out145 = out_145;
assign c_out146 = out_146;
assign c_out147 = out_147;
assign c_out148 = out_148;
assign c_out149 = out_149;
assign c_out150 = out_150;
assign c_out151 = out_151;
assign c_out152 = out_152;
assign c_out153 = out_153;
assign c_out154 = out_154;
assign c_out155 = out_155;
assign c_out156 = out_156;
assign c_out157 = out_157;
assign c_out158 = out_158;
assign c_out159 = out_159;
assign c_out160 = out_160;
assign c_out161 = out_161;
assign c_out162 = out_162;
assign c_out163 = out_163;
assign c_out164 = out_164;
assign c_out165 = out_165;
assign c_out166 = out_166;
assign c_out167 = out_167;
assign c_out168 = out_168;
assign c_out169 = out_169;
assign c_out170 = out_170;
assign c_out171 = out_171;
assign c_out172 = out_172;
assign c_out173 = out_173;
assign c_out174 = out_174;
assign c_out175 = out_175;
assign c_out176 = out_176;
assign c_out177 = out_177;
assign c_out178 = out_178;
assign c_out179 = out_179;
assign c_out180 = out_180;
assign c_out181 = out_181;
assign c_out182 = out_182;
assign c_out183 = out_183;
assign c_out184 = out_184;
assign c_out185 = out_185;
assign c_out186 = out_186;
assign c_out187 = out_187;
assign c_out188 = out_188;
assign c_out189 = out_189;
assign c_out190 = out_190;
assign c_out191 = out_191;
assign c_out192 = out_192;
assign c_out193 = out_193;
assign c_out194 = out_194;
assign c_out195 = out_195;
assign c_out196 = out_196;
assign c_out197 = out_197;
assign c_out198 = out_198;
assign c_out199 = out_199;
assign c_out200 = out_200;
assign c_out201 = out_201;
assign c_out202 = out_202;
assign c_out203 = out_203;
assign c_out204 = out_204;
assign c_out205 = out_205;
assign c_out206 = out_206;
assign c_out207 = out_207;
assign c_out208 = out_208;
assign c_out209 = out_209;
assign c_out210 = out_210;
assign c_out211 = out_211;
assign c_out212 = out_212;
assign c_out213 = out_213;
assign c_out214 = out_214;
assign c_out215 = out_215;
assign c_out216 = out_216;
assign c_out217 = out_217;
assign c_out218 = out_218;
assign c_out219 = out_219;
assign c_out220 = out_220;
assign c_out221 = out_221;
assign c_out222 = out_222;
assign c_out223 = out_223;
assign c_out224 = out_224;
assign c_out225 = out_225;
assign c_out226 = out_226;
assign c_out227 = out_227;
assign c_out228 = out_228;
assign c_out229 = out_229;
assign c_out230 = out_230;
assign c_out231 = out_231;
assign c_out232 = out_232;
assign c_out233 = out_233;
assign c_out234 = out_234;
assign c_out235 = out_235;
assign c_out236 = out_236;
assign c_out237 = out_237;
assign c_out238 = out_238;
assign c_out239 = out_239;
assign c_out240 = out_240;
assign c_out241 = out_241;
assign c_out242 = out_242;
assign c_out243 = out_243;
assign c_out244 = out_244;
assign c_out245 = out_245;
assign c_out246 = out_246;
assign c_out247 = out_247;
assign c_out248 = out_248;
assign c_out249 = out_249;
assign c_out250 = out_250;
assign c_out251 = out_251;
assign c_out252 = out_252;
assign c_out253 = out_253;
assign c_out254 = out_254;
assign c_out255 = out_255;
assign c_out256 = out_256;
assign c_out257 = out_257;
assign c_out258 = out_258;
assign c_out259 = out_259;
assign c_out260 = out_260;
assign c_out261 = out_261;
assign c_out262 = out_262;
assign c_out263 = out_263;
assign c_out264 = out_264;
assign c_out265 = out_265;
assign c_out266 = out_266;
assign c_out267 = out_267;
assign c_out268 = out_268;
assign c_out269 = out_269;
assign c_out270 = out_270;
assign c_out271 = out_271;
assign c_out272 = out_272;
assign c_out273 = out_273;
assign c_out274 = out_274;
assign c_out275 = out_275;
assign c_out276 = out_276;
assign c_out277 = out_277;
assign c_out278 = out_278;
assign c_out279 = out_279;
assign c_out280 = out_280;
assign c_out281 = out_281;
assign c_out282 = out_282;
assign c_out283 = out_283;
assign c_out284 = out_284;
assign c_out285 = out_285;
assign c_out286 = out_286;
assign c_out287 = out_287;
assign c_out288 = out_288;
assign c_out289 = out_289;
assign c_out290 = out_290;
assign c_out291 = out_291;
assign c_out292 = out_292;
assign c_out293 = out_293;
assign c_out294 = out_294;
assign c_out295 = out_295;
assign c_out296 = out_296;
assign c_out297 = out_297;
assign c_out298 = out_298;
assign c_out299 = out_299;
assign c_out300 = out_300;
assign c_out301 = out_301;
assign c_out302 = out_302;
assign c_out303 = out_303;
assign c_out304 = out_304;
assign c_out305 = out_305;
assign c_out306 = out_306;
assign c_out307 = out_307;
assign c_out308 = out_308;
assign c_out309 = out_309;
assign c_out310 = out_310;
assign c_out311 = out_311;
assign c_out312 = out_312;
assign c_out313 = out_313;
assign c_out314 = out_314;
assign c_out315 = out_315;
assign c_out316 = out_316;
assign c_out317 = out_317;
assign c_out318 = out_318;
assign c_out319 = out_319;
assign c_out320 = out_320;
assign c_out321 = out_321;
assign c_out322 = out_322;
assign c_out323 = out_323;
assign c_out324 = out_324;
assign c_out325 = out_325;
assign c_out326 = out_326;
assign c_out327 = out_327;
assign c_out328 = out_328;
assign c_out329 = out_329;
assign c_out330 = out_330;
assign c_out331 = out_331;
assign c_out332 = out_332;
assign c_out333 = out_333;
assign c_out334 = out_334;
assign c_out335 = out_335;
assign c_out336 = out_336;
assign c_out337 = out_337;
assign c_out338 = out_338;
assign c_out339 = out_339;
assign c_out340 = out_340;
assign c_out341 = out_341;
assign c_out342 = out_342;
assign c_out343 = out_343;
assign c_out344 = out_344;
assign c_out345 = out_345;
assign c_out346 = out_346;
assign c_out347 = out_347;
assign c_out348 = out_348;
assign c_out349 = out_349;
assign c_out350 = out_350;
assign c_out351 = out_351;
assign c_out352 = out_352;
assign c_out353 = out_353;
assign c_out354 = out_354;
assign c_out355 = out_355;
assign c_out356 = out_356;
assign c_out357 = out_357;
assign c_out358 = out_358;
assign c_out359 = out_359;
assign c_out360 = out_360;
assign c_out361 = out_361;
assign c_out362 = out_362;
assign c_out363 = out_363;
assign c_out364 = out_364;
assign c_out365 = out_365;
assign c_out366 = out_366;
assign c_out367 = out_367;
assign c_out368 = out_368;
assign c_out369 = out_369;
assign c_out370 = out_370;
assign c_out371 = out_371;
assign c_out372 = out_372;
assign c_out373 = out_373;
assign c_out374 = out_374;
assign c_out375 = out_375;
assign c_out376 = out_376;
assign c_out377 = out_377;
assign c_out378 = out_378;
assign c_out379 = out_379;
assign c_out380 = out_380;
assign c_out381 = out_381;
assign c_out382 = out_382;
assign c_out383 = out_383;
assign c_out384 = out_384;
assign c_out385 = out_385;
assign c_out386 = out_386;
assign c_out387 = out_387;
assign c_out388 = out_388;
assign c_out389 = out_389;
assign c_out390 = out_390;
assign c_out391 = out_391;
assign c_out392 = out_392;
assign c_out393 = out_393;
assign c_out394 = out_394;
assign c_out395 = out_395;
assign c_out396 = out_396;
assign c_out397 = out_397;
assign c_out398 = out_398;
assign c_out399 = out_399;
assign c_out400 = out_400;
assign c_out401 = out_401;
assign c_out402 = out_402;
assign c_out403 = out_403;
assign c_out404 = out_404;
assign c_out405 = out_405;
assign c_out406 = out_406;
assign c_out407 = out_407;
assign c_out408 = out_408;
assign c_out409 = out_409;
assign c_out410 = out_410;
assign c_out411 = out_411;
assign c_out412 = out_412;
assign c_out413 = out_413;
assign c_out414 = out_414;
assign c_out415 = out_415;
assign c_out416 = out_416;
assign c_out417 = out_417;
assign c_out418 = out_418;
assign c_out419 = out_419;
assign c_out420 = out_420;
assign c_out421 = out_421;
assign c_out422 = out_422;
assign c_out423 = out_423;
assign c_out424 = out_424;
assign c_out425 = out_425;
assign c_out426 = out_426;
assign c_out427 = out_427;
assign c_out428 = out_428;
assign c_out429 = out_429;
assign c_out430 = out_430;
assign c_out431 = out_431;
assign c_out432 = out_432;
assign c_out433 = out_433;
assign c_out434 = out_434;
assign c_out435 = out_435;
assign c_out436 = out_436;
assign c_out437 = out_437;
assign c_out438 = out_438;
assign c_out439 = out_439;
assign c_out440 = out_440;
assign c_out441 = out_441;
assign c_out442 = out_442;
assign c_out443 = out_443;
assign c_out444 = out_444;
assign c_out445 = out_445;
assign c_out446 = out_446;
assign c_out447 = out_447;
assign c_out448 = out_448;
assign c_out449 = out_449;
assign c_out450 = out_450;
assign c_out451 = out_451;
assign c_out452 = out_452;
assign c_out453 = out_453;
assign c_out454 = out_454;
assign c_out455 = out_455;
assign c_out456 = out_456;
assign c_out457 = out_457;
assign c_out458 = out_458;
assign c_out459 = out_459;
assign c_out460 = out_460;
assign c_out461 = out_461;
assign c_out462 = out_462;
assign c_out463 = out_463;
assign c_out464 = out_464;
assign c_out465 = out_465;
assign c_out466 = out_466;
assign c_out467 = out_467;
assign c_out468 = out_468;
assign c_out469 = out_469;
assign c_out470 = out_470;
assign c_out471 = out_471;
assign c_out472 = out_472;
assign c_out473 = out_473;
assign c_out474 = out_474;
assign c_out475 = out_475;
assign c_out476 = out_476;
assign c_out477 = out_477;
assign c_out478 = out_478;
assign c_out479 = out_479;
assign c_out480 = out_480;
assign c_out481 = out_481;
assign c_out482 = out_482;
assign c_out483 = out_483;
assign c_out484 = out_484;
assign c_out485 = out_485;
assign c_out486 = out_486;
assign c_out487 = out_487;
assign c_out488 = out_488;
assign c_out489 = out_489;
assign c_out490 = out_490;
assign c_out491 = out_491;
assign c_out492 = out_492;
assign c_out493 = out_493;
assign c_out494 = out_494;
assign c_out495 = out_495;
assign c_out496 = out_496;
assign c_out497 = out_497;
assign c_out498 = out_498;
assign c_out499 = out_499;
assign c_out500 = out_500;
assign c_out501 = out_501;
assign c_out502 = out_502;
assign c_out503 = out_503;
assign c_out504 = out_504;
assign c_out505 = out_505;
assign c_out506 = out_506;
assign c_out507 = out_507;
assign c_out508 = out_508;
assign c_out509 = out_509;
assign c_out510 = out_510;
assign c_out511 = out_511;
assign c_out512 = out_512;
assign c_out513 = out_513;
assign c_out514 = out_514;
assign c_out515 = out_515;
assign c_out516 = out_516;
assign c_out517 = out_517;
assign c_out518 = out_518;
assign c_out519 = out_519;
assign c_out520 = out_520;
assign c_out521 = out_521;
assign c_out522 = out_522;
assign c_out523 = out_523;
assign c_out524 = out_524;
assign c_out525 = out_525;
assign c_out526 = out_526;
assign c_out527 = out_527;
assign c_out528 = out_528;
assign c_out529 = out_529;
assign c_out530 = out_530;
assign c_out531 = out_531;
assign c_out532 = out_532;
assign c_out533 = out_533;
assign c_out534 = out_534;
assign c_out535 = out_535;
assign c_out536 = out_536;
assign c_out537 = out_537;
assign c_out538 = out_538;
assign c_out539 = out_539;
assign c_out540 = out_540;
assign c_out541 = out_541;
assign c_out542 = out_542;
assign c_out543 = out_543;
assign c_out544 = out_544;
assign c_out545 = out_545;
assign c_out546 = out_546;
assign c_out547 = out_547;
assign c_out548 = out_548;
assign c_out549 = out_549;
assign c_out550 = out_550;
assign c_out551 = out_551;
assign c_out552 = out_552;
assign c_out553 = out_553;
assign c_out554 = out_554;
assign c_out555 = out_555;
assign c_out556 = out_556;
assign c_out557 = out_557;
assign c_out558 = out_558;
assign c_out559 = out_559;
assign c_out560 = out_560;
assign c_out561 = out_561;
assign c_out562 = out_562;
assign c_out563 = out_563;
assign c_out564 = out_564;
assign c_out565 = out_565;
assign c_out566 = out_566;
assign c_out567 = out_567;
assign c_out568 = out_568;
assign c_out569 = out_569;
assign c_out570 = out_570;
assign c_out571 = out_571;
assign c_out572 = out_572;
assign c_out573 = out_573;
assign c_out574 = out_574;
assign c_out575 = out_575;
assign c_out576 = out_576;
assign c_out577 = out_577;
assign c_out578 = out_578;
assign c_out579 = out_579;
assign c_out580 = out_580;
assign c_out581 = out_581;
assign c_out582 = out_582;
assign c_out583 = out_583;
assign c_out584 = out_584;
assign c_out585 = out_585;
assign c_out586 = out_586;
assign c_out587 = out_587;
assign c_out588 = out_588;
assign c_out589 = out_589;
assign c_out590 = out_590;
assign c_out591 = out_591;
assign c_out592 = out_592;
assign c_out593 = out_593;
assign c_out594 = out_594;
assign c_out595 = out_595;
assign c_out596 = out_596;
assign c_out597 = out_597;
assign c_out598 = out_598;
assign c_out599 = out_599;
assign c_out600 = out_600;
assign c_out601 = out_601;
assign c_out602 = out_602;
assign c_out603 = out_603;
assign c_out604 = out_604;
assign c_out605 = out_605;
assign c_out606 = out_606;
assign c_out607 = out_607;
assign c_out608 = out_608;
assign c_out609 = out_609;
assign c_out610 = out_610;
assign c_out611 = out_611;
assign c_out612 = out_612;
assign c_out613 = out_613;
assign c_out614 = out_614;
assign c_out615 = out_615;
assign c_out616 = out_616;
assign c_out617 = out_617;
assign c_out618 = out_618;
assign c_out619 = out_619;
assign c_out620 = out_620;
assign c_out621 = out_621;
assign c_out622 = out_622;
assign c_out623 = out_623;
assign c_out624 = out_624;
assign c_out625 = out_625;
assign c_out626 = out_626;
assign c_out627 = out_627;
assign c_out628 = out_628;
assign c_out629 = out_629;
assign c_out630 = out_630;
assign c_out631 = out_631;
assign c_out632 = out_632;
assign c_out633 = out_633;
assign c_out634 = out_634;
assign c_out635 = out_635;
assign c_out636 = out_636;
assign c_out637 = out_637;
assign c_out638 = out_638;
assign c_out639 = out_639;
assign c_out640 = out_640;
assign c_out641 = out_641;
assign c_out642 = out_642;
assign c_out643 = out_643;
assign c_out644 = out_644;
assign c_out645 = out_645;
assign c_out646 = out_646;
assign c_out647 = out_647;
assign c_out648 = out_648;
assign c_out649 = out_649;
assign c_out650 = out_650;
assign c_out651 = out_651;
assign c_out652 = out_652;
assign c_out653 = out_653;
assign c_out654 = out_654;
assign c_out655 = out_655;
assign c_out656 = out_656;
assign c_out657 = out_657;
assign c_out658 = out_658;
assign c_out659 = out_659;
assign c_out660 = out_660;
assign c_out661 = out_661;
assign c_out662 = out_662;
assign c_out663 = out_663;
assign c_out664 = out_664;
assign c_out665 = out_665;
assign c_out666 = out_666;
assign c_out667 = out_667;
assign c_out668 = out_668;
assign c_out669 = out_669;
assign c_out670 = out_670;
assign c_out671 = out_671;
assign c_out672 = out_672;
assign c_out673 = out_673;
assign c_out674 = out_674;
assign c_out675 = out_675;
assign c_out676 = out_676;
assign c_out677 = out_677;
assign c_out678 = out_678;
assign c_out679 = out_679;
assign c_out680 = out_680;
assign c_out681 = out_681;
assign c_out682 = out_682;
assign c_out683 = out_683;
assign c_out684 = out_684;
assign c_out685 = out_685;
assign c_out686 = out_686;
assign c_out687 = out_687;
assign c_out688 = out_688;
assign c_out689 = out_689;
assign c_out690 = out_690;
assign c_out691 = out_691;
assign c_out692 = out_692;
assign c_out693 = out_693;
assign c_out694 = out_694;
assign c_out695 = out_695;
assign c_out696 = out_696;
assign c_out697 = out_697;
assign c_out698 = out_698;
assign c_out699 = out_699;
assign c_out700 = out_700;
assign c_out701 = out_701;
assign c_out702 = out_702;
assign c_out703 = out_703;
assign c_out704 = out_704;
assign c_out705 = out_705;
assign c_out706 = out_706;
assign c_out707 = out_707;
assign c_out708 = out_708;
assign c_out709 = out_709;
assign c_out710 = out_710;
assign c_out711 = out_711;
assign c_out712 = out_712;
assign c_out713 = out_713;
assign c_out714 = out_714;
assign c_out715 = out_715;
assign c_out716 = out_716;
assign c_out717 = out_717;
assign c_out718 = out_718;
assign c_out719 = out_719;
assign c_out720 = out_720;
assign c_out721 = out_721;
assign c_out722 = out_722;
assign c_out723 = out_723;
assign c_out724 = out_724;
assign c_out725 = out_725;
assign c_out726 = out_726;
assign c_out727 = out_727;
assign c_out728 = out_728;
assign c_out729 = out_729;
assign c_out730 = out_730;
assign c_out731 = out_731;
assign c_out732 = out_732;
assign c_out733 = out_733;
assign c_out734 = out_734;
assign c_out735 = out_735;
assign c_out736 = out_736;
assign c_out737 = out_737;
assign c_out738 = out_738;
assign c_out739 = out_739;
assign c_out740 = out_740;
assign c_out741 = out_741;
assign c_out742 = out_742;
assign c_out743 = out_743;
assign c_out744 = out_744;
assign c_out745 = out_745;
assign c_out746 = out_746;
assign c_out747 = out_747;
assign c_out748 = out_748;
assign c_out749 = out_749;
assign c_out750 = out_750;
assign c_out751 = out_751;
assign c_out752 = out_752;
assign c_out753 = out_753;
assign c_out754 = out_754;
assign c_out755 = out_755;
assign c_out756 = out_756;
assign c_out757 = out_757;
assign c_out758 = out_758;
assign c_out759 = out_759;
assign c_out760 = out_760;
assign c_out761 = out_761;
assign c_out762 = out_762;
assign c_out763 = out_763;
assign c_out764 = out_764;
assign c_out765 = out_765;
assign c_out766 = out_766;
assign c_out767 = out_767;
assign c_out768 = out_768;
assign c_out769 = out_769;
assign c_out770 = out_770;
assign c_out771 = out_771;
assign c_out772 = out_772;
assign c_out773 = out_773;
assign c_out774 = out_774;
assign c_out775 = out_775;
assign c_out776 = out_776;
assign c_out777 = out_777;
assign c_out778 = out_778;
assign c_out779 = out_779;
assign c_out780 = out_780;
assign c_out781 = out_781;
assign c_out782 = out_782;
assign c_out783 = out_783;
assign c_out784 = out_784;
assign c_out785 = out_785;
assign c_out786 = out_786;
assign c_out787 = out_787;
assign c_out788 = out_788;
assign c_out789 = out_789;
assign c_out790 = out_790;
assign c_out791 = out_791;
assign c_out792 = out_792;
assign c_out793 = out_793;
assign c_out794 = out_794;
assign c_out795 = out_795;
assign c_out796 = out_796;
assign c_out797 = out_797;
assign c_out798 = out_798;
assign c_out799 = out_799;
assign c_out800 = out_800;
assign c_out801 = out_801;
assign c_out802 = out_802;
assign c_out803 = out_803;
assign c_out804 = out_804;
assign c_out805 = out_805;
assign c_out806 = out_806;
assign c_out807 = out_807;
assign c_out808 = out_808;
assign c_out809 = out_809;
assign c_out810 = out_810;
assign c_out811 = out_811;
assign c_out812 = out_812;
assign c_out813 = out_813;
assign c_out814 = out_814;
assign c_out815 = out_815;
assign c_out816 = out_816;
assign c_out817 = out_817;
assign c_out818 = out_818;
assign c_out819 = out_819;
assign c_out820 = out_820;
assign c_out821 = out_821;
assign c_out822 = out_822;
assign c_out823 = out_823;
assign c_out824 = out_824;
assign c_out825 = out_825;
assign c_out826 = out_826;
assign c_out827 = out_827;
assign c_out828 = out_828;
assign c_out829 = out_829;
assign c_out830 = out_830;
assign c_out831 = out_831;
assign c_out832 = out_832;
assign c_out833 = out_833;
assign c_out834 = out_834;
assign c_out835 = out_835;
assign c_out836 = out_836;
assign c_out837 = out_837;
assign c_out838 = out_838;
assign c_out839 = out_839;
assign c_out840 = out_840;
assign c_out841 = out_841;
assign c_out842 = out_842;
assign c_out843 = out_843;
assign c_out844 = out_844;
assign c_out845 = out_845;
assign c_out846 = out_846;
assign c_out847 = out_847;
assign c_out848 = out_848;
assign c_out849 = out_849;
assign c_out850 = out_850;
assign c_out851 = out_851;
assign c_out852 = out_852;
assign c_out853 = out_853;
assign c_out854 = out_854;
assign c_out855 = out_855;
assign c_out856 = out_856;
assign c_out857 = out_857;
assign c_out858 = out_858;
assign c_out859 = out_859;
assign c_out860 = out_860;
assign c_out861 = out_861;
assign c_out862 = out_862;
assign c_out863 = out_863;
assign c_out864 = out_864;
assign c_out865 = out_865;
assign c_out866 = out_866;
assign c_out867 = out_867;
assign c_out868 = out_868;
assign c_out869 = out_869;
assign c_out870 = out_870;
assign c_out871 = out_871;
assign c_out872 = out_872;
assign c_out873 = out_873;
assign c_out874 = out_874;
assign c_out875 = out_875;
assign c_out876 = out_876;
assign c_out877 = out_877;
assign c_out878 = out_878;
assign c_out879 = out_879;
assign c_out880 = out_880;
assign c_out881 = out_881;
assign c_out882 = out_882;
assign c_out883 = out_883;
assign c_out884 = out_884;
assign c_out885 = out_885;
assign c_out886 = out_886;
assign c_out887 = out_887;
assign c_out888 = out_888;
assign c_out889 = out_889;
assign c_out890 = out_890;
assign c_out891 = out_891;
assign c_out892 = out_892;
assign c_out893 = out_893;
assign c_out894 = out_894;
assign c_out895 = out_895;
assign c_out896 = out_896;
assign c_out897 = out_897;
assign c_out898 = out_898;
assign c_out899 = out_899;
assign c_out900 = out_900;
assign c_out901 = out_901;
assign c_out902 = out_902;
assign c_out903 = out_903;
assign c_out904 = out_904;
assign c_out905 = out_905;
assign c_out906 = out_906;
assign c_out907 = out_907;
assign c_out908 = out_908;
assign c_out909 = out_909;
assign c_out910 = out_910;
assign c_out911 = out_911;
assign c_out912 = out_912;
assign c_out913 = out_913;
assign c_out914 = out_914;
assign c_out915 = out_915;
assign c_out916 = out_916;
assign c_out917 = out_917;
assign c_out918 = out_918;
assign c_out919 = out_919;
assign c_out920 = out_920;
assign c_out921 = out_921;
assign c_out922 = out_922;
assign c_out923 = out_923;
assign c_out924 = out_924;
assign c_out925 = out_925;
assign c_out926 = out_926;
assign c_out927 = out_927;
assign c_out928 = out_928;
assign c_out929 = out_929;
assign c_out930 = out_930;
assign c_out931 = out_931;
assign c_out932 = out_932;
assign c_out933 = out_933;
assign c_out934 = out_934;
assign c_out935 = out_935;
assign c_out936 = out_936;
assign c_out937 = out_937;
assign c_out938 = out_938;
assign c_out939 = out_939;
assign c_out940 = out_940;
assign c_out941 = out_941;
assign c_out942 = out_942;
assign c_out943 = out_943;
assign c_out944 = out_944;
assign c_out945 = out_945;
assign c_out946 = out_946;
assign c_out947 = out_947;
assign c_out948 = out_948;
assign c_out949 = out_949;
assign c_out950 = out_950;
assign c_out951 = out_951;
assign c_out952 = out_952;
assign c_out953 = out_953;
assign c_out954 = out_954;
assign c_out955 = out_955;
assign c_out956 = out_956;
assign c_out957 = out_957;
assign c_out958 = out_958;
assign c_out959 = out_959;
assign c_out960 = out_960;
assign c_out961 = out_961;
assign c_out962 = out_962;
assign c_out963 = out_963;
assign c_out964 = out_964;
assign c_out965 = out_965;
assign c_out966 = out_966;
assign c_out967 = out_967;
assign c_out968 = out_968;
assign c_out969 = out_969;
assign c_out970 = out_970;
assign c_out971 = out_971;
assign c_out972 = out_972;
assign c_out973 = out_973;
assign c_out974 = out_974;
assign c_out975 = out_975;
assign c_out976 = out_976;
assign c_out977 = out_977;
assign c_out978 = out_978;
assign c_out979 = out_979;
assign c_out980 = out_980;
assign c_out981 = out_981;
assign c_out982 = out_982;
assign c_out983 = out_983;
assign c_out984 = out_984;
assign c_out985 = out_985;
assign c_out986 = out_986;
assign c_out987 = out_987;
assign c_out988 = out_988;
assign c_out989 = out_989;
assign c_out990 = out_990;
assign c_out991 = out_991;
assign c_out992 = out_992;
assign c_out993 = out_993;
assign c_out994 = out_994;
assign c_out995 = out_995;
assign c_out996 = out_996;
assign c_out997 = out_997;
assign c_out998 = out_998;
assign c_out999 = out_999;
assign c_out1000 = out_1000;
assign c_out1001 = out_1001;
assign c_out1002 = out_1002;
assign c_out1003 = out_1003;
assign c_out1004 = out_1004;
assign c_out1005 = out_1005;
assign c_out1006 = out_1006;
assign c_out1007 = out_1007;
assign c_out1008 = out_1008;
assign c_out1009 = out_1009;
assign c_out1010 = out_1010;
assign c_out1011 = out_1011;
assign c_out1012 = out_1012;
assign c_out1013 = out_1013;
assign c_out1014 = out_1014;
assign c_out1015 = out_1015;
assign c_out1016 = out_1016;
assign c_out1017 = out_1017;
assign c_out1018 = out_1018;
assign c_out1019 = out_1019;
assign c_out1020 = out_1020;
assign c_out1021 = out_1021;
assign c_out1022 = out_1022;
assign c_out1023 = out_1023;
assign c_out1024 = out_1024;
assign c_out1025 = out_1025;
assign c_out1026 = out_1026;
assign c_out1027 = out_1027;
assign c_out1028 = out_1028;
assign c_out1029 = out_1029;
assign c_out1030 = out_1030;
assign c_out1031 = out_1031;
assign c_out1032 = out_1032;
assign c_out1033 = out_1033;
assign c_out1034 = out_1034;
assign c_out1035 = out_1035;
assign c_out1036 = out_1036;
assign c_out1037 = out_1037;
assign c_out1038 = out_1038;
assign c_out1039 = out_1039;
assign c_out1040 = out_1040;
assign c_out1041 = out_1041;
assign c_out1042 = out_1042;
assign c_out1043 = out_1043;
assign c_out1044 = out_1044;
assign c_out1045 = out_1045;
assign c_out1046 = out_1046;
assign c_out1047 = out_1047;
assign c_out1048 = out_1048;
assign c_out1049 = out_1049;
assign c_out1050 = out_1050;
assign c_out1051 = out_1051;
assign c_out1052 = out_1052;
assign c_out1053 = out_1053;
assign c_out1054 = out_1054;
assign c_out1055 = out_1055;
assign c_out1056 = out_1056;
assign c_out1057 = out_1057;
assign c_out1058 = out_1058;
assign c_out1059 = out_1059;
assign c_out1060 = out_1060;
assign c_out1061 = out_1061;
assign c_out1062 = out_1062;
assign c_out1063 = out_1063;
assign c_out1064 = out_1064;
assign c_out1065 = out_1065;
assign c_out1066 = out_1066;
assign c_out1067 = out_1067;
assign c_out1068 = out_1068;
assign c_out1069 = out_1069;
assign c_out1070 = out_1070;
assign c_out1071 = out_1071;
assign c_out1072 = out_1072;
assign c_out1073 = out_1073;
assign c_out1074 = out_1074;
assign c_out1075 = out_1075;
assign c_out1076 = out_1076;
assign c_out1077 = out_1077;
assign c_out1078 = out_1078;
assign c_out1079 = out_1079;
assign c_out1080 = out_1080;
assign c_out1081 = out_1081;
assign c_out1082 = out_1082;
assign c_out1083 = out_1083;
assign c_out1084 = out_1084;
assign c_out1085 = out_1085;
assign c_out1086 = out_1086;
assign c_out1087 = out_1087;
assign c_out1088 = out_1088;
assign c_out1089 = out_1089;
assign c_out1090 = out_1090;
assign c_out1091 = out_1091;
assign c_out1092 = out_1092;
assign c_out1093 = out_1093;
assign c_out1094 = out_1094;
assign c_out1095 = out_1095;
assign c_out1096 = out_1096;
assign c_out1097 = out_1097;
assign c_out1098 = out_1098;
assign c_out1099 = out_1099;
assign c_out1100 = out_1100;
assign c_out1101 = out_1101;
assign c_out1102 = out_1102;
assign c_out1103 = out_1103;
assign c_out1104 = out_1104;
assign c_out1105 = out_1105;
assign c_out1106 = out_1106;
assign c_out1107 = out_1107;
assign c_out1108 = out_1108;
assign c_out1109 = out_1109;
assign c_out1110 = out_1110;
assign c_out1111 = out_1111;
assign c_out1112 = out_1112;
assign c_out1113 = out_1113;
assign c_out1114 = out_1114;
assign c_out1115 = out_1115;
assign c_out1116 = out_1116;
assign c_out1117 = out_1117;
assign c_out1118 = out_1118;
assign c_out1119 = out_1119;
assign c_out1120 = out_1120;
assign c_out1121 = out_1121;
assign c_out1122 = out_1122;
assign c_out1123 = out_1123;
assign c_out1124 = out_1124;
assign c_out1125 = out_1125;
assign c_out1126 = out_1126;
assign c_out1127 = out_1127;
assign c_out1128 = out_1128;
assign c_out1129 = out_1129;
assign c_out1130 = out_1130;
assign c_out1131 = out_1131;
assign c_out1132 = out_1132;
assign c_out1133 = out_1133;
assign c_out1134 = out_1134;
assign c_out1135 = out_1135;
assign c_out1136 = out_1136;
assign c_out1137 = out_1137;
assign c_out1138 = out_1138;
assign c_out1139 = out_1139;
assign c_out1140 = out_1140;
assign c_out1141 = out_1141;
assign c_out1142 = out_1142;
assign c_out1143 = out_1143;
assign c_out1144 = out_1144;
assign c_out1145 = out_1145;
assign c_out1146 = out_1146;
assign c_out1147 = out_1147;
assign c_out1148 = out_1148;
assign c_out1149 = out_1149;
assign c_out1150 = out_1150;
assign c_out1151 = out_1151;
assign c_out1152 = out_1152;
assign c_out1153 = out_1153;
assign c_out1154 = out_1154;
assign c_out1155 = out_1155;
assign c_out1156 = out_1156;
assign c_out1157 = out_1157;
assign c_out1158 = out_1158;
assign c_out1159 = out_1159;
assign c_out1160 = out_1160;
assign c_out1161 = out_1161;
assign c_out1162 = out_1162;
assign c_out1163 = out_1163;
assign c_out1164 = out_1164;
assign c_out1165 = out_1165;
assign c_out1166 = out_1166;
assign c_out1167 = out_1167;
assign c_out1168 = out_1168;
assign c_out1169 = out_1169;
assign c_out1170 = out_1170;
assign c_out1171 = out_1171;
assign c_out1172 = out_1172;
assign c_out1173 = out_1173;
assign c_out1174 = out_1174;
assign c_out1175 = out_1175;
assign c_out1176 = out_1176;
assign c_out1177 = out_1177;
assign c_out1178 = out_1178;
assign c_out1179 = out_1179;
assign c_out1180 = out_1180;
assign c_out1181 = out_1181;
assign c_out1182 = out_1182;
assign c_out1183 = out_1183;
assign c_out1184 = out_1184;
assign c_out1185 = out_1185;
assign c_out1186 = out_1186;
assign c_out1187 = out_1187;
assign c_out1188 = out_1188;
assign c_out1189 = out_1189;
assign c_out1190 = out_1190;
assign c_out1191 = out_1191;
assign c_out1192 = out_1192;
assign c_out1193 = out_1193;
assign c_out1194 = out_1194;
assign c_out1195 = out_1195;
assign c_out1196 = out_1196;
assign c_out1197 = out_1197;
assign c_out1198 = out_1198;
assign c_out1199 = out_1199;
assign c_out1200 = out_1200;
assign c_out1201 = out_1201;
assign c_out1202 = out_1202;
assign c_out1203 = out_1203;
assign c_out1204 = out_1204;
assign c_out1205 = out_1205;
assign c_out1206 = out_1206;
assign c_out1207 = out_1207;
assign c_out1208 = out_1208;
assign c_out1209 = out_1209;
assign c_out1210 = out_1210;
assign c_out1211 = out_1211;
assign c_out1212 = out_1212;
assign c_out1213 = out_1213;
assign c_out1214 = out_1214;
assign c_out1215 = out_1215;
assign c_out1216 = out_1216;
assign c_out1217 = out_1217;
assign c_out1218 = out_1218;
assign c_out1219 = out_1219;
assign c_out1220 = out_1220;
assign c_out1221 = out_1221;
assign c_out1222 = out_1222;
assign c_out1223 = out_1223;
assign c_out1224 = out_1224;
assign c_out1225 = out_1225;
assign c_out1226 = out_1226;
assign c_out1227 = out_1227;
assign c_out1228 = out_1228;
assign c_out1229 = out_1229;
assign c_out1230 = out_1230;
assign c_out1231 = out_1231;
assign c_out1232 = out_1232;
assign c_out1233 = out_1233;
assign c_out1234 = out_1234;
assign c_out1235 = out_1235;
assign c_out1236 = out_1236;
assign c_out1237 = out_1237;
assign c_out1238 = out_1238;
assign c_out1239 = out_1239;
assign c_out1240 = out_1240;
assign c_out1241 = out_1241;
assign c_out1242 = out_1242;
assign c_out1243 = out_1243;
assign c_out1244 = out_1244;
assign c_out1245 = out_1245;
assign c_out1246 = out_1246;
assign c_out1247 = out_1247;
assign c_out1248 = out_1248;
assign c_out1249 = out_1249;
assign c_out1250 = out_1250;
assign c_out1251 = out_1251;
assign c_out1252 = out_1252;
assign c_out1253 = out_1253;
assign c_out1254 = out_1254;
assign c_out1255 = out_1255;
assign c_out1256 = out_1256;
assign c_out1257 = out_1257;
assign c_out1258 = out_1258;
assign c_out1259 = out_1259;
assign c_out1260 = out_1260;
assign c_out1261 = out_1261;
assign c_out1262 = out_1262;
assign c_out1263 = out_1263;
assign c_out1264 = out_1264;
assign c_out1265 = out_1265;
assign c_out1266 = out_1266;
assign c_out1267 = out_1267;
assign c_out1268 = out_1268;
assign c_out1269 = out_1269;
assign c_out1270 = out_1270;
assign c_out1271 = out_1271;
assign c_out1272 = out_1272;
assign c_out1273 = out_1273;
assign c_out1274 = out_1274;
assign c_out1275 = out_1275;
assign c_out1276 = out_1276;
assign c_out1277 = out_1277;
assign c_out1278 = out_1278;
assign c_out1279 = out_1279;
assign c_out1280 = out_1280;
assign c_out1281 = out_1281;
assign c_out1282 = out_1282;
assign c_out1283 = out_1283;
assign c_out1284 = out_1284;
assign c_out1285 = out_1285;
assign c_out1286 = out_1286;
assign c_out1287 = out_1287;
assign c_out1288 = out_1288;
assign c_out1289 = out_1289;
assign c_out1290 = out_1290;
assign c_out1291 = out_1291;
assign c_out1292 = out_1292;
assign c_out1293 = out_1293;
assign c_out1294 = out_1294;
assign c_out1295 = out_1295;
assign c_out1296 = out_1296;
assign c_out1297 = out_1297;
assign c_out1298 = out_1298;
assign c_out1299 = out_1299;
assign c_out1300 = out_1300;
assign c_out1301 = out_1301;
assign c_out1302 = out_1302;
assign c_out1303 = out_1303;
assign c_out1304 = out_1304;
assign c_out1305 = out_1305;
assign c_out1306 = out_1306;
assign c_out1307 = out_1307;
assign c_out1308 = out_1308;
assign c_out1309 = out_1309;
assign c_out1310 = out_1310;
assign c_out1311 = out_1311;
assign c_out1312 = out_1312;
assign c_out1313 = out_1313;
assign c_out1314 = out_1314;
assign c_out1315 = out_1315;
assign c_out1316 = out_1316;
assign c_out1317 = out_1317;
assign c_out1318 = out_1318;
assign c_out1319 = out_1319;
assign c_out1320 = out_1320;
assign c_out1321 = out_1321;
assign c_out1322 = out_1322;
assign c_out1323 = out_1323;
assign c_out1324 = out_1324;
assign c_out1325 = out_1325;
assign c_out1326 = out_1326;
assign c_out1327 = out_1327;
assign c_out1328 = out_1328;
assign c_out1329 = out_1329;
assign c_out1330 = out_1330;
assign c_out1331 = out_1331;
assign c_out1332 = out_1332;
assign c_out1333 = out_1333;
assign c_out1334 = out_1334;
assign c_out1335 = out_1335;
assign c_out1336 = out_1336;
assign c_out1337 = out_1337;
assign c_out1338 = out_1338;
assign c_out1339 = out_1339;
assign c_out1340 = out_1340;
assign c_out1341 = out_1341;
assign c_out1342 = out_1342;
assign c_out1343 = out_1343;
assign c_out1344 = out_1344;
assign c_out1345 = out_1345;
assign c_out1346 = out_1346;
assign c_out1347 = out_1347;
assign c_out1348 = out_1348;
assign c_out1349 = out_1349;
assign c_out1350 = out_1350;
assign c_out1351 = out_1351;
assign c_out1352 = out_1352;
assign c_out1353 = out_1353;
assign c_out1354 = out_1354;
assign c_out1355 = out_1355;
assign c_out1356 = out_1356;
assign c_out1357 = out_1357;
assign c_out1358 = out_1358;
assign c_out1359 = out_1359;
assign c_out1360 = out_1360;
assign c_out1361 = out_1361;
assign c_out1362 = out_1362;
assign c_out1363 = out_1363;
assign c_out1364 = out_1364;
assign c_out1365 = out_1365;
assign c_out1366 = out_1366;
assign c_out1367 = out_1367;
assign c_out1368 = out_1368;
assign c_out1369 = out_1369;
assign c_out1370 = out_1370;
assign c_out1371 = out_1371;
assign c_out1372 = out_1372;
assign c_out1373 = out_1373;
assign c_out1374 = out_1374;
assign c_out1375 = out_1375;
assign c_out1376 = out_1376;
assign c_out1377 = out_1377;
assign c_out1378 = out_1378;
assign c_out1379 = out_1379;
assign c_out1380 = out_1380;
assign c_out1381 = out_1381;
assign c_out1382 = out_1382;
assign c_out1383 = out_1383;
assign c_out1384 = out_1384;
assign c_out1385 = out_1385;
assign c_out1386 = out_1386;
assign c_out1387 = out_1387;
assign c_out1388 = out_1388;
assign c_out1389 = out_1389;
assign c_out1390 = out_1390;
assign c_out1391 = out_1391;
assign c_out1392 = out_1392;
assign c_out1393 = out_1393;
assign c_out1394 = out_1394;
assign c_out1395 = out_1395;
assign c_out1396 = out_1396;
assign c_out1397 = out_1397;
assign c_out1398 = out_1398;
assign c_out1399 = out_1399;
assign c_out1400 = out_1400;
assign c_out1401 = out_1401;
assign c_out1402 = out_1402;
assign c_out1403 = out_1403;
assign c_out1404 = out_1404;
assign c_out1405 = out_1405;
assign c_out1406 = out_1406;
assign c_out1407 = out_1407;
assign c_out1408 = out_1408;
assign c_out1409 = out_1409;
assign c_out1410 = out_1410;
assign c_out1411 = out_1411;
assign c_out1412 = out_1412;
assign c_out1413 = out_1413;
assign c_out1414 = out_1414;
assign c_out1415 = out_1415;
assign c_out1416 = out_1416;
assign c_out1417 = out_1417;
assign c_out1418 = out_1418;
assign c_out1419 = out_1419;
assign c_out1420 = out_1420;
assign c_out1421 = out_1421;
assign c_out1422 = out_1422;
assign c_out1423 = out_1423;
assign c_out1424 = out_1424;
assign c_out1425 = out_1425;
assign c_out1426 = out_1426;
assign c_out1427 = out_1427;
assign c_out1428 = out_1428;
assign c_out1429 = out_1429;
assign c_out1430 = out_1430;
assign c_out1431 = out_1431;
assign c_out1432 = out_1432;
assign c_out1433 = out_1433;
assign c_out1434 = out_1434;
assign c_out1435 = out_1435;
assign c_out1436 = out_1436;
assign c_out1437 = out_1437;
assign c_out1438 = out_1438;
assign c_out1439 = out_1439;
assign c_out1440 = out_1440;
assign c_out1441 = out_1441;
assign c_out1442 = out_1442;
assign c_out1443 = out_1443;
assign c_out1444 = out_1444;
assign c_out1445 = out_1445;
assign c_out1446 = out_1446;
assign c_out1447 = out_1447;
assign c_out1448 = out_1448;
assign c_out1449 = out_1449;
assign c_out1450 = out_1450;
assign c_out1451 = out_1451;
assign c_out1452 = out_1452;
assign c_out1453 = out_1453;
assign c_out1454 = out_1454;
assign c_out1455 = out_1455;
assign c_out1456 = out_1456;
assign c_out1457 = out_1457;
assign c_out1458 = out_1458;
assign c_out1459 = out_1459;
assign c_out1460 = out_1460;
assign c_out1461 = out_1461;
assign c_out1462 = out_1462;
assign c_out1463 = out_1463;
assign c_out1464 = out_1464;
assign c_out1465 = out_1465;
assign c_out1466 = out_1466;
assign c_out1467 = out_1467;
assign c_out1468 = out_1468;
assign c_out1469 = out_1469;
assign c_out1470 = out_1470;
assign c_out1471 = out_1471;
assign c_out1472 = out_1472;
assign c_out1473 = out_1473;
assign c_out1474 = out_1474;
assign c_out1475 = out_1475;
assign c_out1476 = out_1476;
assign c_out1477 = out_1477;
assign c_out1478 = out_1478;
assign c_out1479 = out_1479;
assign c_out1480 = out_1480;
assign c_out1481 = out_1481;
assign c_out1482 = out_1482;
assign c_out1483 = out_1483;
assign c_out1484 = out_1484;
assign c_out1485 = out_1485;
assign c_out1486 = out_1486;
assign c_out1487 = out_1487;
assign c_out1488 = out_1488;
assign c_out1489 = out_1489;
assign c_out1490 = out_1490;
assign c_out1491 = out_1491;
assign c_out1492 = out_1492;
assign c_out1493 = out_1493;
assign c_out1494 = out_1494;
assign c_out1495 = out_1495;
assign c_out1496 = out_1496;
assign c_out1497 = out_1497;
assign c_out1498 = out_1498;
assign c_out1499 = out_1499;
assign c_out1500 = out_1500;
assign c_out1501 = out_1501;
assign c_out1502 = out_1502;
assign c_out1503 = out_1503;
assign c_out1504 = out_1504;
assign c_out1505 = out_1505;
assign c_out1506 = out_1506;
assign c_out1507 = out_1507;
assign c_out1508 = out_1508;
assign c_out1509 = out_1509;
assign c_out1510 = out_1510;
assign c_out1511 = out_1511;
assign c_out1512 = out_1512;
assign c_out1513 = out_1513;
assign c_out1514 = out_1514;
assign c_out1515 = out_1515;
assign c_out1516 = out_1516;
assign c_out1517 = out_1517;
assign c_out1518 = out_1518;
assign c_out1519 = out_1519;
assign c_out1520 = out_1520;
assign c_out1521 = out_1521;
assign c_out1522 = out_1522;
assign c_out1523 = out_1523;
assign c_out1524 = out_1524;
assign c_out1525 = out_1525;
assign c_out1526 = out_1526;
assign c_out1527 = out_1527;
assign c_out1528 = out_1528;
assign c_out1529 = out_1529;
assign c_out1530 = out_1530;
assign c_out1531 = out_1531;
assign c_out1532 = out_1532;
assign c_out1533 = out_1533;
assign c_out1534 = out_1534;
assign c_out1535 = out_1535;
assign c_out1536 = out_1536;
assign c_out1537 = out_1537;
assign c_out1538 = out_1538;
assign c_out1539 = out_1539;
assign c_out1540 = out_1540;
assign c_out1541 = out_1541;
assign c_out1542 = out_1542;
assign c_out1543 = out_1543;
assign c_out1544 = out_1544;
assign c_out1545 = out_1545;
assign c_out1546 = out_1546;
assign c_out1547 = out_1547;
assign c_out1548 = out_1548;
assign c_out1549 = out_1549;
assign c_out1550 = out_1550;
assign c_out1551 = out_1551;
assign c_out1552 = out_1552;
assign c_out1553 = out_1553;
assign c_out1554 = out_1554;
assign c_out1555 = out_1555;
assign c_out1556 = out_1556;
assign c_out1557 = out_1557;
assign c_out1558 = out_1558;
assign c_out1559 = out_1559;
assign c_out1560 = out_1560;
assign c_out1561 = out_1561;
assign c_out1562 = out_1562;
assign c_out1563 = out_1563;
assign c_out1564 = out_1564;
assign c_out1565 = out_1565;
assign c_out1566 = out_1566;
assign c_out1567 = out_1567;
assign c_out1568 = out_1568;
assign c_out1569 = out_1569;
assign c_out1570 = out_1570;
assign c_out1571 = out_1571;
assign c_out1572 = out_1572;
assign c_out1573 = out_1573;
assign c_out1574 = out_1574;
assign c_out1575 = out_1575;
assign c_out1576 = out_1576;
assign c_out1577 = out_1577;
assign c_out1578 = out_1578;
assign c_out1579 = out_1579;
assign c_out1580 = out_1580;
assign c_out1581 = out_1581;
assign c_out1582 = out_1582;
assign c_out1583 = out_1583;
assign c_out1584 = out_1584;
assign c_out1585 = out_1585;
assign c_out1586 = out_1586;
assign c_out1587 = out_1587;
assign c_out1588 = out_1588;
assign c_out1589 = out_1589;
assign c_out1590 = out_1590;
assign c_out1591 = out_1591;
assign c_out1592 = out_1592;
assign c_out1593 = out_1593;
assign c_out1594 = out_1594;
assign c_out1595 = out_1595;
assign c_out1596 = out_1596;
assign c_out1597 = out_1597;
assign c_out1598 = out_1598;
assign c_out1599 = out_1599;
assign c_out1600 = out_1600;
assign c_out1601 = out_1601;
assign c_out1602 = out_1602;
assign c_out1603 = out_1603;
assign c_out1604 = out_1604;
assign c_out1605 = out_1605;
assign c_out1606 = out_1606;
assign c_out1607 = out_1607;
assign c_out1608 = out_1608;
assign c_out1609 = out_1609;
assign c_out1610 = out_1610;
assign c_out1611 = out_1611;
assign c_out1612 = out_1612;
assign c_out1613 = out_1613;
assign c_out1614 = out_1614;
assign c_out1615 = out_1615;
assign c_out1616 = out_1616;
assign c_out1617 = out_1617;
assign c_out1618 = out_1618;
assign c_out1619 = out_1619;
assign c_out1620 = out_1620;
assign c_out1621 = out_1621;
assign c_out1622 = out_1622;
assign c_out1623 = out_1623;
assign c_out1624 = out_1624;
assign c_out1625 = out_1625;
assign c_out1626 = out_1626;
assign c_out1627 = out_1627;
assign c_out1628 = out_1628;
assign c_out1629 = out_1629;
assign c_out1630 = out_1630;
assign c_out1631 = out_1631;
assign c_out1632 = out_1632;
assign c_out1633 = out_1633;
assign c_out1634 = out_1634;
assign c_out1635 = out_1635;
assign c_out1636 = out_1636;
assign c_out1637 = out_1637;
assign c_out1638 = out_1638;
assign c_out1639 = out_1639;
assign c_out1640 = out_1640;
assign c_out1641 = out_1641;
assign c_out1642 = out_1642;
assign c_out1643 = out_1643;
assign c_out1644 = out_1644;
assign c_out1645 = out_1645;
assign c_out1646 = out_1646;
assign c_out1647 = out_1647;
assign c_out1648 = out_1648;
assign c_out1649 = out_1649;
assign c_out1650 = out_1650;
assign c_out1651 = out_1651;
assign c_out1652 = out_1652;
assign c_out1653 = out_1653;
assign c_out1654 = out_1654;
assign c_out1655 = out_1655;
assign c_out1656 = out_1656;
assign c_out1657 = out_1657;
assign c_out1658 = out_1658;
assign c_out1659 = out_1659;
assign c_out1660 = out_1660;
assign c_out1661 = out_1661;
assign c_out1662 = out_1662;
assign c_out1663 = out_1663;
assign c_out1664 = out_1664;
assign c_out1665 = out_1665;
assign c_out1666 = out_1666;
assign c_out1667 = out_1667;
assign c_out1668 = out_1668;
assign c_out1669 = out_1669;
assign c_out1670 = out_1670;
assign c_out1671 = out_1671;
assign c_out1672 = out_1672;
assign c_out1673 = out_1673;
assign c_out1674 = out_1674;
assign c_out1675 = out_1675;
assign c_out1676 = out_1676;
assign c_out1677 = out_1677;
assign c_out1678 = out_1678;
assign c_out1679 = out_1679;
assign c_out1680 = out_1680;
assign c_out1681 = out_1681;
assign c_out1682 = out_1682;
assign c_out1683 = out_1683;
assign c_out1684 = out_1684;
assign c_out1685 = out_1685;
assign c_out1686 = out_1686;
assign c_out1687 = out_1687;
assign c_out1688 = out_1688;
assign c_out1689 = out_1689;
assign c_out1690 = out_1690;
assign c_out1691 = out_1691;
assign c_out1692 = out_1692;
assign c_out1693 = out_1693;
assign c_out1694 = out_1694;
assign c_out1695 = out_1695;
assign c_out1696 = out_1696;
assign c_out1697 = out_1697;
assign c_out1698 = out_1698;
assign c_out1699 = out_1699;
assign c_out1700 = out_1700;
assign c_out1701 = out_1701;
assign c_out1702 = out_1702;
assign c_out1703 = out_1703;
assign c_out1704 = out_1704;
assign c_out1705 = out_1705;
assign c_out1706 = out_1706;
assign c_out1707 = out_1707;
assign c_out1708 = out_1708;
assign c_out1709 = out_1709;
assign c_out1710 = out_1710;
assign c_out1711 = out_1711;
assign c_out1712 = out_1712;
assign c_out1713 = out_1713;
assign c_out1714 = out_1714;
assign c_out1715 = out_1715;
assign c_out1716 = out_1716;
assign c_out1717 = out_1717;
assign c_out1718 = out_1718;
assign c_out1719 = out_1719;
assign c_out1720 = out_1720;
assign c_out1721 = out_1721;
assign c_out1722 = out_1722;
assign c_out1723 = out_1723;
assign c_out1724 = out_1724;
assign c_out1725 = out_1725;
assign c_out1726 = out_1726;
assign c_out1727 = out_1727;
assign c_out1728 = out_1728;
assign c_out1729 = out_1729;
assign c_out1730 = out_1730;
assign c_out1731 = out_1731;
assign c_out1732 = out_1732;
assign c_out1733 = out_1733;
assign c_out1734 = out_1734;
assign c_out1735 = out_1735;
assign c_out1736 = out_1736;
assign c_out1737 = out_1737;
assign c_out1738 = out_1738;
assign c_out1739 = out_1739;
assign c_out1740 = out_1740;
assign c_out1741 = out_1741;
assign c_out1742 = out_1742;
assign c_out1743 = out_1743;
assign c_out1744 = out_1744;
assign c_out1745 = out_1745;
assign c_out1746 = out_1746;
assign c_out1747 = out_1747;
assign c_out1748 = out_1748;
assign c_out1749 = out_1749;
assign c_out1750 = out_1750;
assign c_out1751 = out_1751;
assign c_out1752 = out_1752;
assign c_out1753 = out_1753;
assign c_out1754 = out_1754;
assign c_out1755 = out_1755;
assign c_out1756 = out_1756;
assign c_out1757 = out_1757;
assign c_out1758 = out_1758;
assign c_out1759 = out_1759;
assign c_out1760 = out_1760;
assign c_out1761 = out_1761;
assign c_out1762 = out_1762;
assign c_out1763 = out_1763;
assign c_out1764 = out_1764;
assign c_out1765 = out_1765;
assign c_out1766 = out_1766;
assign c_out1767 = out_1767;
assign c_out1768 = out_1768;
assign c_out1769 = out_1769;
assign c_out1770 = out_1770;
assign c_out1771 = out_1771;
assign c_out1772 = out_1772;
assign c_out1773 = out_1773;
assign c_out1774 = out_1774;
assign c_out1775 = out_1775;
assign c_out1776 = out_1776;
assign c_out1777 = out_1777;
assign c_out1778 = out_1778;
assign c_out1779 = out_1779;
assign c_out1780 = out_1780;
assign c_out1781 = out_1781;
assign c_out1782 = out_1782;
assign c_out1783 = out_1783;
assign c_out1784 = out_1784;
assign c_out1785 = out_1785;
assign c_out1786 = out_1786;
assign c_out1787 = out_1787;
assign c_out1788 = out_1788;
assign c_out1789 = out_1789;
assign c_out1790 = out_1790;
assign c_out1791 = out_1791;
assign c_out1792 = out_1792;
assign c_out1793 = out_1793;
assign c_out1794 = out_1794;
assign c_out1795 = out_1795;
assign c_out1796 = out_1796;
assign c_out1797 = out_1797;
assign c_out1798 = out_1798;
assign c_out1799 = out_1799;
assign c_out1800 = out_1800;
assign c_out1801 = out_1801;
assign c_out1802 = out_1802;
assign c_out1803 = out_1803;
assign c_out1804 = out_1804;
assign c_out1805 = out_1805;
assign c_out1806 = out_1806;
assign c_out1807 = out_1807;
assign c_out1808 = out_1808;
assign c_out1809 = out_1809;
assign c_out1810 = out_1810;
assign c_out1811 = out_1811;
assign c_out1812 = out_1812;
assign c_out1813 = out_1813;
assign c_out1814 = out_1814;
assign c_out1815 = out_1815;
assign c_out1816 = out_1816;
assign c_out1817 = out_1817;
assign c_out1818 = out_1818;
assign c_out1819 = out_1819;
assign c_out1820 = out_1820;
assign c_out1821 = out_1821;
assign c_out1822 = out_1822;
assign c_out1823 = out_1823;
assign c_out1824 = out_1824;
assign c_out1825 = out_1825;
assign c_out1826 = out_1826;
assign c_out1827 = out_1827;
assign c_out1828 = out_1828;
assign c_out1829 = out_1829;
assign c_out1830 = out_1830;
assign c_out1831 = out_1831;
assign c_out1832 = out_1832;
assign c_out1833 = out_1833;
assign c_out1834 = out_1834;
assign c_out1835 = out_1835;
assign c_out1836 = out_1836;
assign c_out1837 = out_1837;
assign c_out1838 = out_1838;
assign c_out1839 = out_1839;
assign c_out1840 = out_1840;
assign c_out1841 = out_1841;
assign c_out1842 = out_1842;
assign c_out1843 = out_1843;
assign c_out1844 = out_1844;
assign c_out1845 = out_1845;
assign c_out1846 = out_1846;
assign c_out1847 = out_1847;
assign c_out1848 = out_1848;
assign c_out1849 = out_1849;
assign c_out1850 = out_1850;
assign c_out1851 = out_1851;
assign c_out1852 = out_1852;
assign c_out1853 = out_1853;
assign c_out1854 = out_1854;
assign c_out1855 = out_1855;
assign c_out1856 = out_1856;
assign c_out1857 = out_1857;
assign c_out1858 = out_1858;
assign c_out1859 = out_1859;
assign c_out1860 = out_1860;
assign c_out1861 = out_1861;
assign c_out1862 = out_1862;
assign c_out1863 = out_1863;
assign c_out1864 = out_1864;
assign c_out1865 = out_1865;
assign c_out1866 = out_1866;
assign c_out1867 = out_1867;
assign c_out1868 = out_1868;
assign c_out1869 = out_1869;
assign c_out1870 = out_1870;
assign c_out1871 = out_1871;
assign c_out1872 = out_1872;
assign c_out1873 = out_1873;
assign c_out1874 = out_1874;
assign c_out1875 = out_1875;
assign c_out1876 = out_1876;
assign c_out1877 = out_1877;
assign c_out1878 = out_1878;
assign c_out1879 = out_1879;
assign c_out1880 = out_1880;
assign c_out1881 = out_1881;
assign c_out1882 = out_1882;
assign c_out1883 = out_1883;
assign c_out1884 = out_1884;
assign c_out1885 = out_1885;
assign c_out1886 = out_1886;
assign c_out1887 = out_1887;
assign c_out1888 = out_1888;
assign c_out1889 = out_1889;
assign c_out1890 = out_1890;
assign c_out1891 = out_1891;
assign c_out1892 = out_1892;
assign c_out1893 = out_1893;
assign c_out1894 = out_1894;
assign c_out1895 = out_1895;
assign c_out1896 = out_1896;
assign c_out1897 = out_1897;
assign c_out1898 = out_1898;
assign c_out1899 = out_1899;
assign c_out1900 = out_1900;
assign c_out1901 = out_1901;
assign c_out1902 = out_1902;
assign c_out1903 = out_1903;
assign c_out1904 = out_1904;
assign c_out1905 = out_1905;
assign c_out1906 = out_1906;
assign c_out1907 = out_1907;
assign c_out1908 = out_1908;
assign c_out1909 = out_1909;
assign c_out1910 = out_1910;
assign c_out1911 = out_1911;
assign c_out1912 = out_1912;
assign c_out1913 = out_1913;
assign c_out1914 = out_1914;
assign c_out1915 = out_1915;
assign c_out1916 = out_1916;
assign c_out1917 = out_1917;
assign c_out1918 = out_1918;
assign c_out1919 = out_1919;
assign c_out1920 = out_1920;
assign c_out1921 = out_1921;
assign c_out1922 = out_1922;
assign c_out1923 = out_1923;
assign c_out1924 = out_1924;
assign c_out1925 = out_1925;
assign c_out1926 = out_1926;
assign c_out1927 = out_1927;
assign c_out1928 = out_1928;
assign c_out1929 = out_1929;
assign c_out1930 = out_1930;
assign c_out1931 = out_1931;
assign c_out1932 = out_1932;
assign c_out1933 = out_1933;
assign c_out1934 = out_1934;
assign c_out1935 = out_1935;
assign c_out1936 = out_1936;
assign c_out1937 = out_1937;
assign c_out1938 = out_1938;
assign c_out1939 = out_1939;
assign c_out1940 = out_1940;
assign c_out1941 = out_1941;
assign c_out1942 = out_1942;
assign c_out1943 = out_1943;
assign c_out1944 = out_1944;
assign c_out1945 = out_1945;
assign c_out1946 = out_1946;
assign c_out1947 = out_1947;
assign c_out1948 = out_1948;
assign c_out1949 = out_1949;
assign c_out1950 = out_1950;
assign c_out1951 = out_1951;
assign c_out1952 = out_1952;
assign c_out1953 = out_1953;
assign c_out1954 = out_1954;
assign c_out1955 = out_1955;
assign c_out1956 = out_1956;
assign c_out1957 = out_1957;
assign c_out1958 = out_1958;
assign c_out1959 = out_1959;
assign c_out1960 = out_1960;
assign c_out1961 = out_1961;
assign c_out1962 = out_1962;
assign c_out1963 = out_1963;
assign c_out1964 = out_1964;
assign c_out1965 = out_1965;
assign c_out1966 = out_1966;
assign c_out1967 = out_1967;
assign c_out1968 = out_1968;
assign c_out1969 = out_1969;
assign c_out1970 = out_1970;
assign c_out1971 = out_1971;
assign c_out1972 = out_1972;
assign c_out1973 = out_1973;
assign c_out1974 = out_1974;
assign c_out1975 = out_1975;
assign c_out1976 = out_1976;
assign c_out1977 = out_1977;
assign c_out1978 = out_1978;
assign c_out1979 = out_1979;
assign c_out1980 = out_1980;
assign c_out1981 = out_1981;
assign c_out1982 = out_1982;
assign c_out1983 = out_1983;
assign c_out1984 = out_1984;
assign c_out1985 = out_1985;
assign c_out1986 = out_1986;
assign c_out1987 = out_1987;
assign c_out1988 = out_1988;
assign c_out1989 = out_1989;
assign c_out1990 = out_1990;
assign c_out1991 = out_1991;
assign c_out1992 = out_1992;
assign c_out1993 = out_1993;
assign c_out1994 = out_1994;
assign c_out1995 = out_1995;
assign c_out1996 = out_1996;
assign c_out1997 = out_1997;
assign c_out1998 = out_1998;
assign c_out1999 = out_1999;
assign c_out2000 = out_2000;
assign c_out2001 = out_2001;
assign c_out2002 = out_2002;
assign c_out2003 = out_2003;
assign c_out2004 = out_2004;
assign c_out2005 = out_2005;
assign c_out2006 = out_2006;
assign c_out2007 = out_2007;
assign c_out2008 = out_2008;
assign c_out2009 = out_2009;
assign c_out2010 = out_2010;
assign c_out2011 = out_2011;
assign c_out2012 = out_2012;
assign c_out2013 = out_2013;
assign c_out2014 = out_2014;
assign c_out2015 = out_2015;
assign c_out2016 = out_2016;
assign c_out2017 = out_2017;
assign c_out2018 = out_2018;
assign c_out2019 = out_2019;
assign c_out2020 = out_2020;
assign c_out2021 = out_2021;
assign c_out2022 = out_2022;
assign c_out2023 = out_2023;
assign c_out2024 = out_2024;
assign c_out2025 = out_2025;
assign c_out2026 = out_2026;
assign c_out2027 = out_2027;
assign c_out2028 = out_2028;
assign c_out2029 = out_2029;
assign c_out2030 = out_2030;
assign c_out2031 = out_2031;
assign c_out2032 = out_2032;
assign c_out2033 = out_2033;
assign c_out2034 = out_2034;
assign c_out2035 = out_2035;
assign c_out2036 = out_2036;
assign c_out2037 = out_2037;
assign c_out2038 = out_2038;
assign c_out2039 = out_2039;
assign c_out2040 = out_2040;
assign c_out2041 = out_2041;
assign c_out2042 = out_2042;
assign c_out2043 = out_2043;
assign c_out2044 = out_2044;
assign c_out2045 = out_2045;
assign c_out2046 = out_2046;
assign c_out2047 = out_2047;
​


endmodule
