module SA128(clk, rstn, activation, weight, control,c_out0,c_out1,c_out2,c_out3,c_out4,c_out5,c_out6,c_out7,c_out8,c_out9,c_out10,c_out11,c_out12,c_out13,c_out14,c_out15,c_out16,c_out17,c_out18,c_out19,c_out20,c_out21,c_out22,c_out23,c_out24,c_out25,c_out26,c_out27,c_out28,c_out29,c_out30,c_out31,c_out32,c_out33,c_out34,c_out35,c_out36,c_out37,c_out38,c_out39,c_out40,c_out41,c_out42,c_out43,c_out44,c_out45,c_out46,c_out47,c_out48,c_out49,c_out50,c_out51,c_out52,c_out53,c_out54,c_out55,c_out56,c_out57,c_out58,c_out59,c_out60,c_out61,c_out62,c_out63,c_out64,c_out65,c_out66,c_out67,c_out68,c_out69,c_out70,c_out71,c_out72,c_out73,c_out74,c_out75,c_out76,c_out77,c_out78,c_out79,c_out80,c_out81,c_out82,c_out83,c_out84,c_out85,c_out86,c_out87,c_out88,c_out89,c_out90,c_out91,c_out92,c_out93,c_out94,c_out95,c_out96,c_out97,c_out98,c_out99,c_out100,c_out101,c_out102,c_out103,c_out104,c_out105,c_out106,c_out107,c_out108,c_out109,c_out110,c_out111,c_out112,c_out113,c_out114,c_out115,c_out116,c_out117,c_out118,c_out119,c_out120,c_out121,c_out122,c_out123,c_out124,c_out125,c_out126,c_out127,c_out128,c_out129,c_out130,c_out131,c_out132,c_out133,c_out134,c_out135,c_out136,c_out137,c_out138,c_out139,c_out140,c_out141,c_out142,c_out143,c_out144,c_out145,c_out146,c_out147,c_out148,c_out149,c_out150,c_out151,c_out152,c_out153,c_out154,c_out155,c_out156,c_out157,c_out158,c_out159,c_out160,c_out161,c_out162,c_out163,c_out164,c_out165,c_out166,c_out167,c_out168,c_out169,c_out170,c_out171,c_out172,c_out173,c_out174,c_out175,c_out176,c_out177,c_out178,c_out179,c_out180,c_out181,c_out182,c_out183,c_out184,c_out185,c_out186,c_out187,c_out188,c_out189,c_out190,c_out191,c_out192,c_out193,c_out194,c_out195,c_out196,c_out197,c_out198,c_out199,c_out200,c_out201,c_out202,c_out203,c_out204,c_out205,c_out206,c_out207,c_out208,c_out209,c_out210,c_out211,c_out212,c_out213,c_out214,c_out215,c_out216,c_out217,c_out218,c_out219,c_out220,c_out221,c_out222,c_out223,c_out224,c_out225,c_out226,c_out227,c_out228,c_out229,c_out230,c_out231,c_out232,c_out233,c_out234,c_out235,c_out236,c_out237,c_out238,c_out239,c_out240,c_out241,c_out242,c_out243,c_out244,c_out245,c_out246,c_out247,c_out248,c_out249,c_out250,c_out251,c_out252,c_out253,c_out254,c_out255,c_out256, c_out257, c_out258, c_out259, c_out260, c_out261, c_out262, c_out263, c_out264, c_out265, c_out266, c_out267, c_out268, c_out269, c_out270, c_out271, c_out272, c_out273,  c_out274, c_out275, c_out276, c_out277, c_out278, c_out279, c_out280, c_out281, c_out282, c_out283, c_out284,  c_out285, c_out286, c_out287, c_out288, c_out289, c_out290, c_out291, c_out292, c_out293, c_out294, c_out295, c_out296, c_out297, c_out298, c_out299, c_out300, c_out301, c_out302, c_out303, c_out304, c_out305, c_out306,c_out307, c_out308,  c_out309, c_out310, c_out311, c_out312, c_out313, c_out314, c_out315, c_out316, c_out317, c_out318, c_out319, c_out320, c_out321, c_out322, c_out323, c_out324, c_out325, c_out326, c_out327, c_out328, c_out329, c_out330, c_out331, c_out332, c_out333, c_out334, c_out335, c_out336, c_out337, c_out338, c_out339, c_out340, c_out341, c_out342, c_out343, c_out344, c_out345, c_out346, c_out347, c_out348, c_out349, c_out350, c_out351, c_out352, c_out353, c_out354, c_out355, c_out356, c_out357, c_out358, c_out359,c_out360,c_out361, c_out362, c_out363, c_out364, c_out365, c_out366, c_out367, c_out368, c_out369, c_out370, c_out371, c_out372, c_out373, c_out374, c_out375, c_out376, c_out377, c_out378, c_out379, c_out380, c_out381, c_out382, c_out383, c_out384, c_out385, c_out386, c_out387, c_out388, c_out389, c_out390, c_out391, c_out392, c_out393, c_out394, c_out395, c_out396, c_out397, c_out398, c_out399, c_out400, c_out401, c_out402, c_out403, c_out404, c_out405, c_out406, c_out407, c_out408, c_out409, c_out410, c_out411, c_out412, c_out413, c_out414, c_out415, c_out416, c_out417, c_out418, c_out419, c_out420, c_out421, c_out422, c_out423, c_out424, c_out425, c_out426, c_out427, c_out428, c_out429, c_out430, c_out431, c_out432, c_out433, c_out434, c_out435, c_out436, c_out437, c_out438, c_out439, c_out440, c_out441, c_out442, c_out443, c_out444, c_out445, c_out446, c_out447, c_out448, c_out449, c_out450, c_out451, c_out452, c_out453, c_out454, c_out455, c_out456, c_out457, c_out458, c_out459, c_out460, c_out461, c_out462, c_out463, c_out464, c_out465, c_out466, c_out467, c_out468, c_out469, c_out470, c_out471, c_out472, c_out473, c_out474, c_out475, c_out476, c_out477, c_out478, c_out479, c_out480, c_out481, c_out482, c_out483, c_out484, c_out485, c_out486, c_out487, c_out488, c_out489, c_out490, c_out491, c_out492, c_out493, c_out494, c_out495, c_out496, c_out497, c_out498, c_out499, c_out500, c_out501, c_out502, c_out503, c_out504, c_out505, c_out506, c_out507, c_out508, c_out509, c_out510, c_out511, out_act,out_weight);
parameter WIDTH = 8;
parameter C_WIDTH = 32;

input clk,rstn;
input [128*WIDTH-1:0] activation;
input [128*WIDTH-1:0] weight;
input control;
output [32*C_WIDTH-1:0] c_out0;
output [32*C_WIDTH-1:0] c_out1;
output [32*C_WIDTH-1:0] c_out2;
output [32*C_WIDTH-1:0] c_out3;
output [32*C_WIDTH-1:0] c_out4;
output [32*C_WIDTH-1:0] c_out5;
output [32*C_WIDTH-1:0] c_out6;
output [32*C_WIDTH-1:0] c_out7;
output [32*C_WIDTH-1:0] c_out8;
output [32*C_WIDTH-1:0] c_out9;
output [32*C_WIDTH-1:0] c_out10;
output [32*C_WIDTH-1:0] c_out11;
output [32*C_WIDTH-1:0] c_out12;
output [32*C_WIDTH-1:0] c_out13;
output [32*C_WIDTH-1:0] c_out14;
output [32*C_WIDTH-1:0] c_out15;
output [32*C_WIDTH-1:0] c_out16;
output [32*C_WIDTH-1:0] c_out17;
output [32*C_WIDTH-1:0] c_out18;
output [32*C_WIDTH-1:0] c_out19;
output [32*C_WIDTH-1:0] c_out20;
output [32*C_WIDTH-1:0] c_out21;
output [32*C_WIDTH-1:0] c_out22;
output [32*C_WIDTH-1:0] c_out23;
output [32*C_WIDTH-1:0] c_out24;
output [32*C_WIDTH-1:0] c_out25;
output [32*C_WIDTH-1:0] c_out26;
output [32*C_WIDTH-1:0] c_out27;
output [32*C_WIDTH-1:0] c_out28;
output [32*C_WIDTH-1:0] c_out29;
output [32*C_WIDTH-1:0] c_out30;
output [32*C_WIDTH-1:0] c_out31;
output [32*C_WIDTH-1:0] c_out32;
output [32*C_WIDTH-1:0] c_out33;
output [32*C_WIDTH-1:0] c_out34;
output [32*C_WIDTH-1:0] c_out35;
output [32*C_WIDTH-1:0] c_out36;
output [32*C_WIDTH-1:0] c_out37;
output [32*C_WIDTH-1:0] c_out38;
output [32*C_WIDTH-1:0] c_out39;
output [32*C_WIDTH-1:0] c_out40;
output [32*C_WIDTH-1:0] c_out41;
output [32*C_WIDTH-1:0] c_out42;
output [32*C_WIDTH-1:0] c_out43;
output [32*C_WIDTH-1:0] c_out44;
output [32*C_WIDTH-1:0] c_out45;
output [32*C_WIDTH-1:0] c_out46;
output [32*C_WIDTH-1:0] c_out47;
output [32*C_WIDTH-1:0] c_out48;
output [32*C_WIDTH-1:0] c_out49;
output [32*C_WIDTH-1:0] c_out50;
output [32*C_WIDTH-1:0] c_out51;
output [32*C_WIDTH-1:0] c_out52;
output [32*C_WIDTH-1:0] c_out53;
output [32*C_WIDTH-1:0] c_out54;
output [32*C_WIDTH-1:0] c_out55;
output [32*C_WIDTH-1:0] c_out56;
output [32*C_WIDTH-1:0] c_out57;
output [32*C_WIDTH-1:0] c_out58;
output [32*C_WIDTH-1:0] c_out59;
output [32*C_WIDTH-1:0] c_out60;
output [32*C_WIDTH-1:0] c_out61;
output [32*C_WIDTH-1:0] c_out62;
output [32*C_WIDTH-1:0] c_out63;
output [32*C_WIDTH-1:0] c_out64;
output [32*C_WIDTH-1:0] c_out65;
output [32*C_WIDTH-1:0] c_out66;
output [32*C_WIDTH-1:0] c_out67;
output [32*C_WIDTH-1:0] c_out68;
output [32*C_WIDTH-1:0] c_out69;
output [32*C_WIDTH-1:0] c_out70;
output [32*C_WIDTH-1:0] c_out71;
output [32*C_WIDTH-1:0] c_out72;
output [32*C_WIDTH-1:0] c_out73;
output [32*C_WIDTH-1:0] c_out74;
output [32*C_WIDTH-1:0] c_out75;
output [32*C_WIDTH-1:0] c_out76;
output [32*C_WIDTH-1:0] c_out77;
output [32*C_WIDTH-1:0] c_out78;
output [32*C_WIDTH-1:0] c_out79;
output [32*C_WIDTH-1:0] c_out80;
output [32*C_WIDTH-1:0] c_out81;
output [32*C_WIDTH-1:0] c_out82;
output [32*C_WIDTH-1:0] c_out83;
output [32*C_WIDTH-1:0] c_out84;
output [32*C_WIDTH-1:0] c_out85;
output [32*C_WIDTH-1:0] c_out86;
output [32*C_WIDTH-1:0] c_out87;
output [32*C_WIDTH-1:0] c_out88;
output [32*C_WIDTH-1:0] c_out89;
output [32*C_WIDTH-1:0] c_out90;
output [32*C_WIDTH-1:0] c_out91;
output [32*C_WIDTH-1:0] c_out92;
output [32*C_WIDTH-1:0] c_out93;
output [32*C_WIDTH-1:0] c_out94;
output [32*C_WIDTH-1:0] c_out95;
output [32*C_WIDTH-1:0] c_out96;
output [32*C_WIDTH-1:0] c_out97;
output [32*C_WIDTH-1:0] c_out98;
output [32*C_WIDTH-1:0] c_out99;
output [32*C_WIDTH-1:0] c_out100;
output [32*C_WIDTH-1:0] c_out101;
output [32*C_WIDTH-1:0] c_out102;
output [32*C_WIDTH-1:0] c_out103;
output [32*C_WIDTH-1:0] c_out104;
output [32*C_WIDTH-1:0] c_out105;
output [32*C_WIDTH-1:0] c_out106;
output [32*C_WIDTH-1:0] c_out107;
output [32*C_WIDTH-1:0] c_out108;
output [32*C_WIDTH-1:0] c_out109;
output [32*C_WIDTH-1:0] c_out110;
output [32*C_WIDTH-1:0] c_out111;
output [32*C_WIDTH-1:0] c_out112;
output [32*C_WIDTH-1:0] c_out113;
output [32*C_WIDTH-1:0] c_out114;
output [32*C_WIDTH-1:0] c_out115;
output [32*C_WIDTH-1:0] c_out116;
output [32*C_WIDTH-1:0] c_out117;
output [32*C_WIDTH-1:0] c_out118;
output [32*C_WIDTH-1:0] c_out119;
output [32*C_WIDTH-1:0] c_out120;
output [32*C_WIDTH-1:0] c_out121;
output [32*C_WIDTH-1:0] c_out122;
output [32*C_WIDTH-1:0] c_out123;
output [32*C_WIDTH-1:0] c_out124;
output [32*C_WIDTH-1:0] c_out125;
output [32*C_WIDTH-1:0] c_out126;
output [32*C_WIDTH-1:0] c_out127;
output [32*C_WIDTH-1:0] c_out128;
output [32*C_WIDTH-1:0] c_out129;
output [32*C_WIDTH-1:0] c_out130;
output [32*C_WIDTH-1:0] c_out131;
output [32*C_WIDTH-1:0] c_out132;
output [32*C_WIDTH-1:0] c_out133;
output [32*C_WIDTH-1:0] c_out134;
output [32*C_WIDTH-1:0] c_out135;
output [32*C_WIDTH-1:0] c_out136;
output [32*C_WIDTH-1:0] c_out137;
output [32*C_WIDTH-1:0] c_out138;
output [32*C_WIDTH-1:0] c_out139;
output [32*C_WIDTH-1:0] c_out140;
output [32*C_WIDTH-1:0] c_out141;
output [32*C_WIDTH-1:0] c_out142;
output [32*C_WIDTH-1:0] c_out143;
output [32*C_WIDTH-1:0] c_out144;
output [32*C_WIDTH-1:0] c_out145;
output [32*C_WIDTH-1:0] c_out146;
output [32*C_WIDTH-1:0] c_out147;
output [32*C_WIDTH-1:0] c_out148;
output [32*C_WIDTH-1:0] c_out149;
output [32*C_WIDTH-1:0] c_out150;
output [32*C_WIDTH-1:0] c_out151;
output [32*C_WIDTH-1:0] c_out152;
output [32*C_WIDTH-1:0] c_out153;
output [32*C_WIDTH-1:0] c_out154;
output [32*C_WIDTH-1:0] c_out155;
output [32*C_WIDTH-1:0] c_out156;
output [32*C_WIDTH-1:0] c_out157;
output [32*C_WIDTH-1:0] c_out158;
output [32*C_WIDTH-1:0] c_out159;
output [32*C_WIDTH-1:0] c_out160;
output [32*C_WIDTH-1:0] c_out161;
output [32*C_WIDTH-1:0] c_out162;
output [32*C_WIDTH-1:0] c_out163;
output [32*C_WIDTH-1:0] c_out164;
output [32*C_WIDTH-1:0] c_out165;
output [32*C_WIDTH-1:0] c_out166;
output [32*C_WIDTH-1:0] c_out167;
output [32*C_WIDTH-1:0] c_out168;
output [32*C_WIDTH-1:0] c_out169;
output [32*C_WIDTH-1:0] c_out170;
output [32*C_WIDTH-1:0] c_out171;
output [32*C_WIDTH-1:0] c_out172;
output [32*C_WIDTH-1:0] c_out173;
output [32*C_WIDTH-1:0] c_out174;
output [32*C_WIDTH-1:0] c_out175;
output [32*C_WIDTH-1:0] c_out176;
output [32*C_WIDTH-1:0] c_out177;
output [32*C_WIDTH-1:0] c_out178;
output [32*C_WIDTH-1:0] c_out179;
output [32*C_WIDTH-1:0] c_out180;
output [32*C_WIDTH-1:0] c_out181;
output [32*C_WIDTH-1:0] c_out182;
output [32*C_WIDTH-1:0] c_out183;
output [32*C_WIDTH-1:0] c_out184;
output [32*C_WIDTH-1:0] c_out185;
output [32*C_WIDTH-1:0] c_out186;
output [32*C_WIDTH-1:0] c_out187;
output [32*C_WIDTH-1:0] c_out188;
output [32*C_WIDTH-1:0] c_out189;
output [32*C_WIDTH-1:0] c_out190;
output [32*C_WIDTH-1:0] c_out191;
output [32*C_WIDTH-1:0] c_out192;
output [32*C_WIDTH-1:0] c_out193;
output [32*C_WIDTH-1:0] c_out194;
output [32*C_WIDTH-1:0] c_out195;
output [32*C_WIDTH-1:0] c_out196;
output [32*C_WIDTH-1:0] c_out197;
output [32*C_WIDTH-1:0] c_out198;
output [32*C_WIDTH-1:0] c_out199;
output [32*C_WIDTH-1:0] c_out200;
output [32*C_WIDTH-1:0] c_out201;
output [32*C_WIDTH-1:0] c_out202;
output [32*C_WIDTH-1:0] c_out203;
output [32*C_WIDTH-1:0] c_out204;
output [32*C_WIDTH-1:0] c_out205;
output [32*C_WIDTH-1:0] c_out206;
output [32*C_WIDTH-1:0] c_out207;
output [32*C_WIDTH-1:0] c_out208;
output [32*C_WIDTH-1:0] c_out209;
output [32*C_WIDTH-1:0] c_out210;
output [32*C_WIDTH-1:0] c_out211;
output [32*C_WIDTH-1:0] c_out212;
output [32*C_WIDTH-1:0] c_out213;
output [32*C_WIDTH-1:0] c_out214;
output [32*C_WIDTH-1:0] c_out215;
output [32*C_WIDTH-1:0] c_out216;
output [32*C_WIDTH-1:0] c_out217;
output [32*C_WIDTH-1:0] c_out218;
output [32*C_WIDTH-1:0] c_out219;
output [32*C_WIDTH-1:0] c_out220;
output [32*C_WIDTH-1:0] c_out221;
output [32*C_WIDTH-1:0] c_out222;
output [32*C_WIDTH-1:0] c_out223;
output [32*C_WIDTH-1:0] c_out224;
output [32*C_WIDTH-1:0] c_out225;
output [32*C_WIDTH-1:0] c_out226;
output [32*C_WIDTH-1:0] c_out227;
output [32*C_WIDTH-1:0] c_out228;
output [32*C_WIDTH-1:0] c_out229;
output [32*C_WIDTH-1:0] c_out230;
output [32*C_WIDTH-1:0] c_out231;
output [32*C_WIDTH-1:0] c_out232;
output [32*C_WIDTH-1:0] c_out233;
output [32*C_WIDTH-1:0] c_out234;
output [32*C_WIDTH-1:0] c_out235;
output [32*C_WIDTH-1:0] c_out236;
output [32*C_WIDTH-1:0] c_out237;
output [32*C_WIDTH-1:0] c_out238;
output [32*C_WIDTH-1:0] c_out239;
output [32*C_WIDTH-1:0] c_out240;
output [32*C_WIDTH-1:0] c_out241;
output [32*C_WIDTH-1:0] c_out242;
output [32*C_WIDTH-1:0] c_out243;
output [32*C_WIDTH-1:0] c_out244;
output [32*C_WIDTH-1:0] c_out245;
output [32*C_WIDTH-1:0] c_out246;
output [32*C_WIDTH-1:0] c_out247;
output [32*C_WIDTH-1:0] c_out248;
output [32*C_WIDTH-1:0] c_out249;
output [32*C_WIDTH-1:0] c_out250;
output [32*C_WIDTH-1:0] c_out251;
output [32*C_WIDTH-1:0] c_out252;
output [32*C_WIDTH-1:0] c_out253;
output [32*C_WIDTH-1:0] c_out254;
output [32*C_WIDTH-1:0] c_out255;
output [32*C_WIDTH-1:0] c_out256;
output [32*C_WIDTH-1:0] c_out257;
output [32*C_WIDTH-1:0] c_out258;
output [32*C_WIDTH-1:0] c_out259;
output [32*C_WIDTH-1:0] c_out260;
output [32*C_WIDTH-1:0] c_out261;
output [32*C_WIDTH-1:0] c_out262;
output [32*C_WIDTH-1:0] c_out263;
output [32*C_WIDTH-1:0] c_out264;
output [32*C_WIDTH-1:0] c_out265;
output [32*C_WIDTH-1:0] c_out266;
output [32*C_WIDTH-1:0] c_out267;
output [32*C_WIDTH-1:0] c_out268;
output [32*C_WIDTH-1:0] c_out269;
output [32*C_WIDTH-1:0] c_out270;
output [32*C_WIDTH-1:0] c_out271;
output [32*C_WIDTH-1:0] c_out272;
output [32*C_WIDTH-1:0] c_out273;
output [32*C_WIDTH-1:0] c_out274;
output [32*C_WIDTH-1:0] c_out275;
output [32*C_WIDTH-1:0] c_out276;
output [32*C_WIDTH-1:0] c_out277;
output [32*C_WIDTH-1:0] c_out278;
output [32*C_WIDTH-1:0] c_out279;
output [32*C_WIDTH-1:0] c_out280;
output [32*C_WIDTH-1:0] c_out281;
output [32*C_WIDTH-1:0] c_out282;
output [32*C_WIDTH-1:0] c_out283;
output [32*C_WIDTH-1:0] c_out284;
output [32*C_WIDTH-1:0] c_out285;
output [32*C_WIDTH-1:0] c_out286;
output [32*C_WIDTH-1:0] c_out287;
output [32*C_WIDTH-1:0] c_out288;
output [32*C_WIDTH-1:0] c_out289;
output [32*C_WIDTH-1:0] c_out290;
output [32*C_WIDTH-1:0] c_out291;
output [32*C_WIDTH-1:0] c_out292;
output [32*C_WIDTH-1:0] c_out293;
output [32*C_WIDTH-1:0] c_out294;
output [32*C_WIDTH-1:0] c_out295;
output [32*C_WIDTH-1:0] c_out296;
output [32*C_WIDTH-1:0] c_out297;
output [32*C_WIDTH-1:0] c_out298;
output [32*C_WIDTH-1:0] c_out299;
output [32*C_WIDTH-1:0] c_out300;
output [32*C_WIDTH-1:0] c_out301;
output [32*C_WIDTH-1:0] c_out302;
output [32*C_WIDTH-1:0] c_out303;
output [32*C_WIDTH-1:0] c_out304;
output [32*C_WIDTH-1:0] c_out305;
output [32*C_WIDTH-1:0] c_out306;
output [32*C_WIDTH-1:0] c_out307;
output [32*C_WIDTH-1:0] c_out308;
output [32*C_WIDTH-1:0] c_out309;
output [32*C_WIDTH-1:0] c_out310;
output [32*C_WIDTH-1:0] c_out311;
output [32*C_WIDTH-1:0] c_out312;
output [32*C_WIDTH-1:0] c_out313;
output [32*C_WIDTH-1:0] c_out314;
output [32*C_WIDTH-1:0] c_out315;
output [32*C_WIDTH-1:0] c_out316;
output [32*C_WIDTH-1:0] c_out317;
output [32*C_WIDTH-1:0] c_out318;
output [32*C_WIDTH-1:0] c_out319;
output [32*C_WIDTH-1:0] c_out320;
output [32*C_WIDTH-1:0] c_out321;
output [32*C_WIDTH-1:0] c_out322;
output [32*C_WIDTH-1:0] c_out323;
output [32*C_WIDTH-1:0] c_out324;
output [32*C_WIDTH-1:0] c_out325;
output [32*C_WIDTH-1:0] c_out326;
output [32*C_WIDTH-1:0] c_out327;
output [32*C_WIDTH-1:0] c_out328;
output [32*C_WIDTH-1:0] c_out329;
output [32*C_WIDTH-1:0] c_out330;
output [32*C_WIDTH-1:0] c_out331;
output [32*C_WIDTH-1:0] c_out332;
output [32*C_WIDTH-1:0] c_out333;
output [32*C_WIDTH-1:0] c_out334;
output [32*C_WIDTH-1:0] c_out335;
output [32*C_WIDTH-1:0] c_out336;
output [32*C_WIDTH-1:0] c_out337;
output [32*C_WIDTH-1:0] c_out338;
output [32*C_WIDTH-1:0] c_out339;
output [32*C_WIDTH-1:0] c_out340;
output [32*C_WIDTH-1:0] c_out341;
output [32*C_WIDTH-1:0] c_out342;
output [32*C_WIDTH-1:0] c_out343;
output [32*C_WIDTH-1:0] c_out344;
output [32*C_WIDTH-1:0] c_out345;
output [32*C_WIDTH-1:0] c_out346;
output [32*C_WIDTH-1:0] c_out347;
output [32*C_WIDTH-1:0] c_out348;
output [32*C_WIDTH-1:0] c_out349;
output [32*C_WIDTH-1:0] c_out350;
output [32*C_WIDTH-1:0] c_out351;
output [32*C_WIDTH-1:0] c_out352;
output [32*C_WIDTH-1:0] c_out353;
output [32*C_WIDTH-1:0] c_out354;
output [32*C_WIDTH-1:0] c_out355;
output [32*C_WIDTH-1:0] c_out356;
output [32*C_WIDTH-1:0] c_out357;
output [32*C_WIDTH-1:0] c_out358;
output [32*C_WIDTH-1:0] c_out359;
output [32*C_WIDTH-1:0] c_out360;
output [32*C_WIDTH-1:0] c_out361;
output [32*C_WIDTH-1:0] c_out362;
output [32*C_WIDTH-1:0] c_out363;
output [32*C_WIDTH-1:0] c_out364;
output [32*C_WIDTH-1:0] c_out365;
output [32*C_WIDTH-1:0] c_out366;
output [32*C_WIDTH-1:0] c_out367;
output [32*C_WIDTH-1:0] c_out368;
output [32*C_WIDTH-1:0] c_out369;
output [32*C_WIDTH-1:0] c_out370;
output [32*C_WIDTH-1:0] c_out371;
output [32*C_WIDTH-1:0] c_out372;
output [32*C_WIDTH-1:0] c_out373;
output [32*C_WIDTH-1:0] c_out374;
output [32*C_WIDTH-1:0] c_out375;
output [32*C_WIDTH-1:0] c_out376;
output [32*C_WIDTH-1:0] c_out377;
output [32*C_WIDTH-1:0] c_out378;
output [32*C_WIDTH-1:0] c_out379;
output [32*C_WIDTH-1:0] c_out380;
output [32*C_WIDTH-1:0] c_out381;
output [32*C_WIDTH-1:0] c_out382;
output [32*C_WIDTH-1:0] c_out383;
output [32*C_WIDTH-1:0] c_out384;
output [32*C_WIDTH-1:0] c_out385;
output [32*C_WIDTH-1:0] c_out386;
output [32*C_WIDTH-1:0] c_out387;
output [32*C_WIDTH-1:0] c_out388;
output [32*C_WIDTH-1:0] c_out389;
output [32*C_WIDTH-1:0] c_out390;
output [32*C_WIDTH-1:0] c_out391;
output [32*C_WIDTH-1:0] c_out392;
output [32*C_WIDTH-1:0] c_out393;
output [32*C_WIDTH-1:0] c_out394;
output [32*C_WIDTH-1:0] c_out395;
output [32*C_WIDTH-1:0] c_out396;
output [32*C_WIDTH-1:0] c_out397;
output [32*C_WIDTH-1:0] c_out398;
output [32*C_WIDTH-1:0] c_out399;
output [32*C_WIDTH-1:0] c_out400;
output [32*C_WIDTH-1:0] c_out401;
output [32*C_WIDTH-1:0] c_out402;
output [32*C_WIDTH-1:0] c_out403;
output [32*C_WIDTH-1:0] c_out404;
output [32*C_WIDTH-1:0] c_out405;
output [32*C_WIDTH-1:0] c_out406;
output [32*C_WIDTH-1:0] c_out407;
output [32*C_WIDTH-1:0] c_out408;
output [32*C_WIDTH-1:0] c_out409;
output [32*C_WIDTH-1:0] c_out410;
output [32*C_WIDTH-1:0] c_out411;
output [32*C_WIDTH-1:0] c_out412;
output [32*C_WIDTH-1:0] c_out413;
output [32*C_WIDTH-1:0] c_out414;
output [32*C_WIDTH-1:0] c_out415;
output [32*C_WIDTH-1:0] c_out416;
output [32*C_WIDTH-1:0] c_out417;
output [32*C_WIDTH-1:0] c_out418;
output [32*C_WIDTH-1:0] c_out419;
output [32*C_WIDTH-1:0] c_out420;
output [32*C_WIDTH-1:0] c_out421;
output [32*C_WIDTH-1:0] c_out422;
output [32*C_WIDTH-1:0] c_out423;
output [32*C_WIDTH-1:0] c_out424;
output [32*C_WIDTH-1:0] c_out425;
output [32*C_WIDTH-1:0] c_out426;
output [32*C_WIDTH-1:0] c_out427;
output [32*C_WIDTH-1:0] c_out428;
output [32*C_WIDTH-1:0] c_out429;
output [32*C_WIDTH-1:0] c_out430;
output [32*C_WIDTH-1:0] c_out431;
output [32*C_WIDTH-1:0] c_out432;
output [32*C_WIDTH-1:0] c_out433;
output [32*C_WIDTH-1:0] c_out434;
output [32*C_WIDTH-1:0] c_out435;
output [32*C_WIDTH-1:0] c_out436;
output [32*C_WIDTH-1:0] c_out437;
output [32*C_WIDTH-1:0] c_out438;
output [32*C_WIDTH-1:0] c_out439;
output [32*C_WIDTH-1:0] c_out440;
output [32*C_WIDTH-1:0] c_out441;
output [32*C_WIDTH-1:0] c_out442;
output [32*C_WIDTH-1:0] c_out443;
output [32*C_WIDTH-1:0] c_out444;
output [32*C_WIDTH-1:0] c_out445;
output [32*C_WIDTH-1:0] c_out446;
output [32*C_WIDTH-1:0] c_out447;
output [32*C_WIDTH-1:0] c_out448;
output [32*C_WIDTH-1:0] c_out449;
output [32*C_WIDTH-1:0] c_out450;
output [32*C_WIDTH-1:0] c_out451;
output [32*C_WIDTH-1:0] c_out452;
output [32*C_WIDTH-1:0] c_out453;
output [32*C_WIDTH-1:0] c_out454;
output [32*C_WIDTH-1:0] c_out455;
output [32*C_WIDTH-1:0] c_out456;
output [32*C_WIDTH-1:0] c_out457;
output [32*C_WIDTH-1:0] c_out458;
output [32*C_WIDTH-1:0] c_out459;
output [32*C_WIDTH-1:0] c_out460;
output [32*C_WIDTH-1:0] c_out461;
output [32*C_WIDTH-1:0] c_out462;
output [32*C_WIDTH-1:0] c_out463;
output [32*C_WIDTH-1:0] c_out464;
output [32*C_WIDTH-1:0] c_out465;
output [32*C_WIDTH-1:0] c_out466;
output [32*C_WIDTH-1:0] c_out467;
output [32*C_WIDTH-1:0] c_out468;
output [32*C_WIDTH-1:0] c_out469;
output [32*C_WIDTH-1:0] c_out470;
output [32*C_WIDTH-1:0] c_out471;
output [32*C_WIDTH-1:0] c_out472;
output [32*C_WIDTH-1:0] c_out473;
output [32*C_WIDTH-1:0] c_out474;
output [32*C_WIDTH-1:0] c_out475;
output [32*C_WIDTH-1:0] c_out476;
output [32*C_WIDTH-1:0] c_out477;
output [32*C_WIDTH-1:0] c_out478;
output [32*C_WIDTH-1:0] c_out479;
output [32*C_WIDTH-1:0] c_out480;
output [32*C_WIDTH-1:0] c_out481;
output [32*C_WIDTH-1:0] c_out482;
output [32*C_WIDTH-1:0] c_out483;
output [32*C_WIDTH-1:0] c_out484;
output [32*C_WIDTH-1:0] c_out485;
output [32*C_WIDTH-1:0] c_out486;
output [32*C_WIDTH-1:0] c_out487;
output [32*C_WIDTH-1:0] c_out488;
output [32*C_WIDTH-1:0] c_out489;
output [32*C_WIDTH-1:0] c_out490;
output [32*C_WIDTH-1:0] c_out491;
output [32*C_WIDTH-1:0] c_out492;
output [32*C_WIDTH-1:0] c_out493;
output [32*C_WIDTH-1:0] c_out494;
output [32*C_WIDTH-1:0] c_out495;
output [32*C_WIDTH-1:0] c_out496;
output [32*C_WIDTH-1:0] c_out497;
output [32*C_WIDTH-1:0] c_out498;
output [32*C_WIDTH-1:0] c_out499;
output [32*C_WIDTH-1:0] c_out500;
output [32*C_WIDTH-1:0] c_out501;
output [32*C_WIDTH-1:0] c_out502;
output [32*C_WIDTH-1:0] c_out503;
output [32*C_WIDTH-1:0] c_out504;
output [32*C_WIDTH-1:0] c_out505;
output [32*C_WIDTH-1:0] c_out506;
output [32*C_WIDTH-1:0] c_out507;
output [32*C_WIDTH-1:0] c_out508;
output [32*C_WIDTH-1:0] c_out509;
output [32*C_WIDTH-1:0] c_out510;
output [32*C_WIDTH-1:0] c_out511;

output [128*WIDTH-1:0] out_act;
output [128*WIDTH-1:0] out_weight;


wire [64*WIDTH-1:0] act_0;
wire [64*WIDTH-1:0] act_1;
wire [64*WIDTH-1:0] weight_0;
wire [64*WIDTH-1:0] weight_1;

wire [64*WIDTH-1:0] outact_0;
wire [64*WIDTH-1:0] outact_1;
wire [64*WIDTH-1:0] outweight_0;
wire [64*WIDTH-1:0] outweight_1;

wire [64*WIDTH-1:0] act0_1;
wire [64*WIDTH-1:0] act2_3;
wire [64*WIDTH-1:0] weight0_2;
wire [64*WIDTH-1:0] weight1_3;
wire [32*C_WIDTH-1:0] out_0;
wire [32*C_WIDTH-1:0] out_1;
wire [32*C_WIDTH-1:0] out_2;
wire [32*C_WIDTH-1:0] out_3;
wire [32*C_WIDTH-1:0] out_4;
wire [32*C_WIDTH-1:0] out_5;
wire [32*C_WIDTH-1:0] out_6;
wire [32*C_WIDTH-1:0] out_7;
wire [32*C_WIDTH-1:0] out_8;
wire [32*C_WIDTH-1:0] out_9;
wire [32*C_WIDTH-1:0] out_10;
wire [32*C_WIDTH-1:0] out_11;
wire [32*C_WIDTH-1:0] out_12;
wire [32*C_WIDTH-1:0] out_13;
wire [32*C_WIDTH-1:0] out_14;
wire [32*C_WIDTH-1:0] out_15;
wire [32*C_WIDTH-1:0] out_16;
wire [32*C_WIDTH-1:0] out_17;
wire [32*C_WIDTH-1:0] out_18;
wire [32*C_WIDTH-1:0] out_19;
wire [32*C_WIDTH-1:0] out_20;
wire [32*C_WIDTH-1:0] out_21;
wire [32*C_WIDTH-1:0] out_22;
wire [32*C_WIDTH-1:0] out_23;
wire [32*C_WIDTH-1:0] out_24;
wire [32*C_WIDTH-1:0] out_25;
wire [32*C_WIDTH-1:0] out_26;
wire [32*C_WIDTH-1:0] out_27;
wire [32*C_WIDTH-1:0] out_28;
wire [32*C_WIDTH-1:0] out_29;
wire [32*C_WIDTH-1:0] out_30;
wire [32*C_WIDTH-1:0] out_31;
wire [32*C_WIDTH-1:0] out_32;
wire [32*C_WIDTH-1:0] out_33;
wire [32*C_WIDTH-1:0] out_34;
wire [32*C_WIDTH-1:0] out_35;
wire [32*C_WIDTH-1:0] out_36;
wire [32*C_WIDTH-1:0] out_37;
wire [32*C_WIDTH-1:0] out_38;
wire [32*C_WIDTH-1:0] out_39;
wire [32*C_WIDTH-1:0] out_40;
wire [32*C_WIDTH-1:0] out_41;
wire [32*C_WIDTH-1:0] out_42;
wire [32*C_WIDTH-1:0] out_43;
wire [32*C_WIDTH-1:0] out_44;
wire [32*C_WIDTH-1:0] out_45;
wire [32*C_WIDTH-1:0] out_46;
wire [32*C_WIDTH-1:0] out_47;
wire [32*C_WIDTH-1:0] out_48;
wire [32*C_WIDTH-1:0] out_49;
wire [32*C_WIDTH-1:0] out_50;
wire [32*C_WIDTH-1:0] out_51;
wire [32*C_WIDTH-1:0] out_52;
wire [32*C_WIDTH-1:0] out_53;
wire [32*C_WIDTH-1:0] out_54;
wire [32*C_WIDTH-1:0] out_55;
wire [32*C_WIDTH-1:0] out_56;
wire [32*C_WIDTH-1:0] out_57;
wire [32*C_WIDTH-1:0] out_58;
wire [32*C_WIDTH-1:0] out_59;
wire [32*C_WIDTH-1:0] out_60;
wire [32*C_WIDTH-1:0] out_61;
wire [32*C_WIDTH-1:0] out_62;
wire [32*C_WIDTH-1:0] out_63;
wire [32*C_WIDTH-1:0] out_64;
wire [32*C_WIDTH-1:0] out_65;
wire [32*C_WIDTH-1:0] out_66;
wire [32*C_WIDTH-1:0] out_67;
wire [32*C_WIDTH-1:0] out_68;
wire [32*C_WIDTH-1:0] out_69;
wire [32*C_WIDTH-1:0] out_70;
wire [32*C_WIDTH-1:0] out_71;
wire [32*C_WIDTH-1:0] out_72;
wire [32*C_WIDTH-1:0] out_73;
wire [32*C_WIDTH-1:0] out_74;
wire [32*C_WIDTH-1:0] out_75;
wire [32*C_WIDTH-1:0] out_76;
wire [32*C_WIDTH-1:0] out_77;
wire [32*C_WIDTH-1:0] out_78;
wire [32*C_WIDTH-1:0] out_79;
wire [32*C_WIDTH-1:0] out_80;
wire [32*C_WIDTH-1:0] out_81;
wire [32*C_WIDTH-1:0] out_82;
wire [32*C_WIDTH-1:0] out_83;
wire [32*C_WIDTH-1:0] out_84;
wire [32*C_WIDTH-1:0] out_85;
wire [32*C_WIDTH-1:0] out_86;
wire [32*C_WIDTH-1:0] out_87;
wire [32*C_WIDTH-1:0] out_88;
wire [32*C_WIDTH-1:0] out_89;
wire [32*C_WIDTH-1:0] out_90;
wire [32*C_WIDTH-1:0] out_91;
wire [32*C_WIDTH-1:0] out_92;
wire [32*C_WIDTH-1:0] out_93;
wire [32*C_WIDTH-1:0] out_94;
wire [32*C_WIDTH-1:0] out_95;
wire [32*C_WIDTH-1:0] out_96;
wire [32*C_WIDTH-1:0] out_97;
wire [32*C_WIDTH-1:0] out_98;
wire [32*C_WIDTH-1:0] out_99;
wire [32*C_WIDTH-1:0] out_100;
wire [32*C_WIDTH-1:0] out_101;
wire [32*C_WIDTH-1:0] out_102;
wire [32*C_WIDTH-1:0] out_103;
wire [32*C_WIDTH-1:0] out_104;
wire [32*C_WIDTH-1:0] out_105;
wire [32*C_WIDTH-1:0] out_106;
wire [32*C_WIDTH-1:0] out_107;
wire [32*C_WIDTH-1:0] out_108;
wire [32*C_WIDTH-1:0] out_109;
wire [32*C_WIDTH-1:0] out_110;
wire [32*C_WIDTH-1:0] out_111;
wire [32*C_WIDTH-1:0] out_112;
wire [32*C_WIDTH-1:0] out_113;
wire [32*C_WIDTH-1:0] out_114;
wire [32*C_WIDTH-1:0] out_115;
wire [32*C_WIDTH-1:0] out_116;
wire [32*C_WIDTH-1:0] out_117;
wire [32*C_WIDTH-1:0] out_118;
wire [32*C_WIDTH-1:0] out_119;
wire [32*C_WIDTH-1:0] out_120;
wire [32*C_WIDTH-1:0] out_121;
wire [32*C_WIDTH-1:0] out_122;
wire [32*C_WIDTH-1:0] out_123;
wire [32*C_WIDTH-1:0] out_124;
wire [32*C_WIDTH-1:0] out_125;
wire [32*C_WIDTH-1:0] out_126;
wire [32*C_WIDTH-1:0] out_127;
wire [32*C_WIDTH-1:0] out_128;
wire [32*C_WIDTH-1:0] out_129;
wire [32*C_WIDTH-1:0] out_130;
wire [32*C_WIDTH-1:0] out_131;
wire [32*C_WIDTH-1:0] out_132;
wire [32*C_WIDTH-1:0] out_133;
wire [32*C_WIDTH-1:0] out_134;
wire [32*C_WIDTH-1:0] out_135;
wire [32*C_WIDTH-1:0] out_136;
wire [32*C_WIDTH-1:0] out_137;
wire [32*C_WIDTH-1:0] out_138;
wire [32*C_WIDTH-1:0] out_139;
wire [32*C_WIDTH-1:0] out_140;
wire [32*C_WIDTH-1:0] out_141;
wire [32*C_WIDTH-1:0] out_142;
wire [32*C_WIDTH-1:0] out_143;
wire [32*C_WIDTH-1:0] out_144;
wire [32*C_WIDTH-1:0] out_145;
wire [32*C_WIDTH-1:0] out_146;
wire [32*C_WIDTH-1:0] out_147;
wire [32*C_WIDTH-1:0] out_148;
wire [32*C_WIDTH-1:0] out_149;
wire [32*C_WIDTH-1:0] out_150;
wire [32*C_WIDTH-1:0] out_151;
wire [32*C_WIDTH-1:0] out_152;
wire [32*C_WIDTH-1:0] out_153;
wire [32*C_WIDTH-1:0] out_154;
wire [32*C_WIDTH-1:0] out_155;
wire [32*C_WIDTH-1:0] out_156;
wire [32*C_WIDTH-1:0] out_157;
wire [32*C_WIDTH-1:0] out_158;
wire [32*C_WIDTH-1:0] out_159;
wire [32*C_WIDTH-1:0] out_160;
wire [32*C_WIDTH-1:0] out_161;
wire [32*C_WIDTH-1:0] out_162;
wire [32*C_WIDTH-1:0] out_163;
wire [32*C_WIDTH-1:0] out_164;
wire [32*C_WIDTH-1:0] out_165;
wire [32*C_WIDTH-1:0] out_166;
wire [32*C_WIDTH-1:0] out_167;
wire [32*C_WIDTH-1:0] out_168;
wire [32*C_WIDTH-1:0] out_169;
wire [32*C_WIDTH-1:0] out_170;
wire [32*C_WIDTH-1:0] out_171;
wire [32*C_WIDTH-1:0] out_172;
wire [32*C_WIDTH-1:0] out_173;
wire [32*C_WIDTH-1:0] out_174;
wire [32*C_WIDTH-1:0] out_175;
wire [32*C_WIDTH-1:0] out_176;
wire [32*C_WIDTH-1:0] out_177;
wire [32*C_WIDTH-1:0] out_178;
wire [32*C_WIDTH-1:0] out_179;
wire [32*C_WIDTH-1:0] out_180;
wire [32*C_WIDTH-1:0] out_181;
wire [32*C_WIDTH-1:0] out_182;
wire [32*C_WIDTH-1:0] out_183;
wire [32*C_WIDTH-1:0] out_184;
wire [32*C_WIDTH-1:0] out_185;
wire [32*C_WIDTH-1:0] out_186;
wire [32*C_WIDTH-1:0] out_187;
wire [32*C_WIDTH-1:0] out_188;
wire [32*C_WIDTH-1:0] out_189;
wire [32*C_WIDTH-1:0] out_190;
wire [32*C_WIDTH-1:0] out_191;
wire [32*C_WIDTH-1:0] out_192;
wire [32*C_WIDTH-1:0] out_193;
wire [32*C_WIDTH-1:0] out_194;
wire [32*C_WIDTH-1:0] out_195;
wire [32*C_WIDTH-1:0] out_196;
wire [32*C_WIDTH-1:0] out_197;
wire [32*C_WIDTH-1:0] out_198;
wire [32*C_WIDTH-1:0] out_199;
wire [32*C_WIDTH-1:0] out_200;
wire [32*C_WIDTH-1:0] out_201;
wire [32*C_WIDTH-1:0] out_202;
wire [32*C_WIDTH-1:0] out_203;
wire [32*C_WIDTH-1:0] out_204;
wire [32*C_WIDTH-1:0] out_205;
wire [32*C_WIDTH-1:0] out_206;
wire [32*C_WIDTH-1:0] out_207;
wire [32*C_WIDTH-1:0] out_208;
wire [32*C_WIDTH-1:0] out_209;
wire [32*C_WIDTH-1:0] out_210;
wire [32*C_WIDTH-1:0] out_211;
wire [32*C_WIDTH-1:0] out_212;
wire [32*C_WIDTH-1:0] out_213;
wire [32*C_WIDTH-1:0] out_214;
wire [32*C_WIDTH-1:0] out_215;
wire [32*C_WIDTH-1:0] out_216;
wire [32*C_WIDTH-1:0] out_217;
wire [32*C_WIDTH-1:0] out_218;
wire [32*C_WIDTH-1:0] out_219;
wire [32*C_WIDTH-1:0] out_220;
wire [32*C_WIDTH-1:0] out_221;
wire [32*C_WIDTH-1:0] out_222;
wire [32*C_WIDTH-1:0] out_223;
wire [32*C_WIDTH-1:0] out_224;
wire [32*C_WIDTH-1:0] out_225;
wire [32*C_WIDTH-1:0] out_226;
wire [32*C_WIDTH-1:0] out_227;
wire [32*C_WIDTH-1:0] out_228;
wire [32*C_WIDTH-1:0] out_229;
wire [32*C_WIDTH-1:0] out_230;
wire [32*C_WIDTH-1:0] out_231;
wire [32*C_WIDTH-1:0] out_232;
wire [32*C_WIDTH-1:0] out_233;
wire [32*C_WIDTH-1:0] out_234;
wire [32*C_WIDTH-1:0] out_235;
wire [32*C_WIDTH-1:0] out_236;
wire [32*C_WIDTH-1:0] out_237;
wire [32*C_WIDTH-1:0] out_238;
wire [32*C_WIDTH-1:0] out_239;
wire [32*C_WIDTH-1:0] out_240;
wire [32*C_WIDTH-1:0] out_241;
wire [32*C_WIDTH-1:0] out_242;
wire [32*C_WIDTH-1:0] out_243;
wire [32*C_WIDTH-1:0] out_244;
wire [32*C_WIDTH-1:0] out_245;
wire [32*C_WIDTH-1:0] out_246;
wire [32*C_WIDTH-1:0] out_247;
wire [32*C_WIDTH-1:0] out_248;
wire [32*C_WIDTH-1:0] out_249;
wire [32*C_WIDTH-1:0] out_250;
wire [32*C_WIDTH-1:0] out_251;
wire [32*C_WIDTH-1:0] out_252;
wire [32*C_WIDTH-1:0] out_253;
wire [32*C_WIDTH-1:0] out_254;
wire [32*C_WIDTH-1:0] out_255;
wire [32*C_WIDTH-1:0] out_256;
wire [32*C_WIDTH-1:0] out_257;
wire [32*C_WIDTH-1:0] out_258;
wire [32*C_WIDTH-1:0] out_259;
wire [32*C_WIDTH-1:0] out_260;
wire [32*C_WIDTH-1:0] out_261;
wire [32*C_WIDTH-1:0] out_262;
wire [32*C_WIDTH-1:0] out_263;
wire [32*C_WIDTH-1:0] out_264;
wire [32*C_WIDTH-1:0] out_265;
wire [32*C_WIDTH-1:0] out_266;
wire [32*C_WIDTH-1:0] out_267;
wire [32*C_WIDTH-1:0] out_268;
wire [32*C_WIDTH-1:0] out_269;
wire [32*C_WIDTH-1:0] out_270;
wire [32*C_WIDTH-1:0] out_271;
wire [32*C_WIDTH-1:0] out_272;
wire [32*C_WIDTH-1:0] out_273;
wire [32*C_WIDTH-1:0] out_274;
wire [32*C_WIDTH-1:0] out_275;
wire [32*C_WIDTH-1:0] out_276;
wire [32*C_WIDTH-1:0] out_277;
wire [32*C_WIDTH-1:0] out_278;
wire [32*C_WIDTH-1:0] out_279;
wire [32*C_WIDTH-1:0] out_280;
wire [32*C_WIDTH-1:0] out_281;
wire [32*C_WIDTH-1:0] out_282;
wire [32*C_WIDTH-1:0] out_283;
wire [32*C_WIDTH-1:0] out_284;
wire [32*C_WIDTH-1:0] out_285;
wire [32*C_WIDTH-1:0] out_286;
wire [32*C_WIDTH-1:0] out_287;
wire [32*C_WIDTH-1:0] out_288;
wire [32*C_WIDTH-1:0] out_289;
wire [32*C_WIDTH-1:0] out_290;
wire [32*C_WIDTH-1:0] out_291;
wire [32*C_WIDTH-1:0] out_292;
wire [32*C_WIDTH-1:0] out_293;
wire [32*C_WIDTH-1:0] out_294;
wire [32*C_WIDTH-1:0] out_295;
wire [32*C_WIDTH-1:0] out_296;
wire [32*C_WIDTH-1:0] out_297;
wire [32*C_WIDTH-1:0] out_298;
wire [32*C_WIDTH-1:0] out_299;
wire [32*C_WIDTH-1:0] out_300;
wire [32*C_WIDTH-1:0] out_301;
wire [32*C_WIDTH-1:0] out_302;
wire [32*C_WIDTH-1:0] out_303;
wire [32*C_WIDTH-1:0] out_304;
wire [32*C_WIDTH-1:0] out_305;
wire [32*C_WIDTH-1:0] out_306;
wire [32*C_WIDTH-1:0] out_307;
wire [32*C_WIDTH-1:0] out_308;
wire [32*C_WIDTH-1:0] out_309;
wire [32*C_WIDTH-1:0] out_310;
wire [32*C_WIDTH-1:0] out_311;
wire [32*C_WIDTH-1:0] out_312;
wire [32*C_WIDTH-1:0] out_313;
wire [32*C_WIDTH-1:0] out_314;
wire [32*C_WIDTH-1:0] out_315;
wire [32*C_WIDTH-1:0] out_316;
wire [32*C_WIDTH-1:0] out_317;
wire [32*C_WIDTH-1:0] out_318;
wire [32*C_WIDTH-1:0] out_319;
wire [32*C_WIDTH-1:0] out_320;
wire [32*C_WIDTH-1:0] out_321;
wire [32*C_WIDTH-1:0] out_322;
wire [32*C_WIDTH-1:0] out_323;
wire [32*C_WIDTH-1:0] out_324;
wire [32*C_WIDTH-1:0] out_325;
wire [32*C_WIDTH-1:0] out_326;
wire [32*C_WIDTH-1:0] out_327;
wire [32*C_WIDTH-1:0] out_328;
wire [32*C_WIDTH-1:0] out_329;
wire [32*C_WIDTH-1:0] out_330;
wire [32*C_WIDTH-1:0] out_331;
wire [32*C_WIDTH-1:0] out_332;
wire [32*C_WIDTH-1:0] out_333;
wire [32*C_WIDTH-1:0] out_334;
wire [32*C_WIDTH-1:0] out_335;
wire [32*C_WIDTH-1:0] out_336;
wire [32*C_WIDTH-1:0] out_337;
wire [32*C_WIDTH-1:0] out_338;
wire [32*C_WIDTH-1:0] out_339;
wire [32*C_WIDTH-1:0] out_340;
wire [32*C_WIDTH-1:0] out_341;
wire [32*C_WIDTH-1:0] out_342;
wire [32*C_WIDTH-1:0] out_343;
wire [32*C_WIDTH-1:0] out_344;
wire [32*C_WIDTH-1:0] out_345;
wire [32*C_WIDTH-1:0] out_346;
wire [32*C_WIDTH-1:0] out_347;
wire [32*C_WIDTH-1:0] out_348;
wire [32*C_WIDTH-1:0] out_349;
wire [32*C_WIDTH-1:0] out_350;
wire [32*C_WIDTH-1:0] out_351;
wire [32*C_WIDTH-1:0] out_352;
wire [32*C_WIDTH-1:0] out_353;
wire [32*C_WIDTH-1:0] out_354;
wire [32*C_WIDTH-1:0] out_355;
wire [32*C_WIDTH-1:0] out_356;
wire [32*C_WIDTH-1:0] out_357;
wire [32*C_WIDTH-1:0] out_358;
wire [32*C_WIDTH-1:0] out_359;
wire [32*C_WIDTH-1:0] out_360;
wire [32*C_WIDTH-1:0] out_361;
wire [32*C_WIDTH-1:0] out_362;
wire [32*C_WIDTH-1:0] out_363;
wire [32*C_WIDTH-1:0] out_364;
wire [32*C_WIDTH-1:0] out_365;
wire [32*C_WIDTH-1:0] out_366;
wire [32*C_WIDTH-1:0] out_367;
wire [32*C_WIDTH-1:0] out_368;
wire [32*C_WIDTH-1:0] out_369;
wire [32*C_WIDTH-1:0] out_370;
wire [32*C_WIDTH-1:0] out_371;
wire [32*C_WIDTH-1:0] out_372;
wire [32*C_WIDTH-1:0] out_373;
wire [32*C_WIDTH-1:0] out_374;
wire [32*C_WIDTH-1:0] out_375;
wire [32*C_WIDTH-1:0] out_376;
wire [32*C_WIDTH-1:0] out_377;
wire [32*C_WIDTH-1:0] out_378;
wire [32*C_WIDTH-1:0] out_379;
wire [32*C_WIDTH-1:0] out_380;
wire [32*C_WIDTH-1:0] out_381;
wire [32*C_WIDTH-1:0] out_382;
wire [32*C_WIDTH-1:0] out_383;
wire [32*C_WIDTH-1:0] out_384;
wire [32*C_WIDTH-1:0] out_385;
wire [32*C_WIDTH-1:0] out_386;
wire [32*C_WIDTH-1:0] out_387;
wire [32*C_WIDTH-1:0] out_388;
wire [32*C_WIDTH-1:0] out_389;
wire [32*C_WIDTH-1:0] out_390;
wire [32*C_WIDTH-1:0] out_391;
wire [32*C_WIDTH-1:0] out_392;
wire [32*C_WIDTH-1:0] out_393;
wire [32*C_WIDTH-1:0] out_394;
wire [32*C_WIDTH-1:0] out_395;
wire [32*C_WIDTH-1:0] out_396;
wire [32*C_WIDTH-1:0] out_397;
wire [32*C_WIDTH-1:0] out_398;
wire [32*C_WIDTH-1:0] out_399;
wire [32*C_WIDTH-1:0] out_400;
wire [32*C_WIDTH-1:0] out_401;
wire [32*C_WIDTH-1:0] out_402;
wire [32*C_WIDTH-1:0] out_403;
wire [32*C_WIDTH-1:0] out_404;
wire [32*C_WIDTH-1:0] out_405;
wire [32*C_WIDTH-1:0] out_406;
wire [32*C_WIDTH-1:0] out_407;
wire [32*C_WIDTH-1:0] out_408;
wire [32*C_WIDTH-1:0] out_409;
wire [32*C_WIDTH-1:0] out_410;
wire [32*C_WIDTH-1:0] out_411;
wire [32*C_WIDTH-1:0] out_412;
wire [32*C_WIDTH-1:0] out_413;
wire [32*C_WIDTH-1:0] out_414;
wire [32*C_WIDTH-1:0] out_415;
wire [32*C_WIDTH-1:0] out_416;
wire [32*C_WIDTH-1:0] out_417;
wire [32*C_WIDTH-1:0] out_418;
wire [32*C_WIDTH-1:0] out_419;
wire [32*C_WIDTH-1:0] out_420;
wire [32*C_WIDTH-1:0] out_421;
wire [32*C_WIDTH-1:0] out_422;
wire [32*C_WIDTH-1:0] out_423;
wire [32*C_WIDTH-1:0] out_424;
wire [32*C_WIDTH-1:0] out_425;
wire [32*C_WIDTH-1:0] out_426;
wire [32*C_WIDTH-1:0] out_427;
wire [32*C_WIDTH-1:0] out_428;
wire [32*C_WIDTH-1:0] out_429;
wire [32*C_WIDTH-1:0] out_430;
wire [32*C_WIDTH-1:0] out_431;
wire [32*C_WIDTH-1:0] out_432;
wire [32*C_WIDTH-1:0] out_433;
wire [32*C_WIDTH-1:0] out_434;
wire [32*C_WIDTH-1:0] out_435;
wire [32*C_WIDTH-1:0] out_436;
wire [32*C_WIDTH-1:0] out_437;
wire [32*C_WIDTH-1:0] out_438;
wire [32*C_WIDTH-1:0] out_439;
wire [32*C_WIDTH-1:0] out_440;
wire [32*C_WIDTH-1:0] out_441;
wire [32*C_WIDTH-1:0] out_442;
wire [32*C_WIDTH-1:0] out_443;
wire [32*C_WIDTH-1:0] out_444;
wire [32*C_WIDTH-1:0] out_445;
wire [32*C_WIDTH-1:0] out_446;
wire [32*C_WIDTH-1:0] out_447;
wire [32*C_WIDTH-1:0] out_448;
wire [32*C_WIDTH-1:0] out_449;
wire [32*C_WIDTH-1:0] out_450;
wire [32*C_WIDTH-1:0] out_451;
wire [32*C_WIDTH-1:0] out_452;
wire [32*C_WIDTH-1:0] out_453;
wire [32*C_WIDTH-1:0] out_454;
wire [32*C_WIDTH-1:0] out_455;
wire [32*C_WIDTH-1:0] out_456;
wire [32*C_WIDTH-1:0] out_457;
wire [32*C_WIDTH-1:0] out_458;
wire [32*C_WIDTH-1:0] out_459;
wire [32*C_WIDTH-1:0] out_460;
wire [32*C_WIDTH-1:0] out_461;
wire [32*C_WIDTH-1:0] out_462;
wire [32*C_WIDTH-1:0] out_463;
wire [32*C_WIDTH-1:0] out_464;
wire [32*C_WIDTH-1:0] out_465;
wire [32*C_WIDTH-1:0] out_466;
wire [32*C_WIDTH-1:0] out_467;
wire [32*C_WIDTH-1:0] out_468;
wire [32*C_WIDTH-1:0] out_469;
wire [32*C_WIDTH-1:0] out_470;
wire [32*C_WIDTH-1:0] out_471;
wire [32*C_WIDTH-1:0] out_472;
wire [32*C_WIDTH-1:0] out_473;
wire [32*C_WIDTH-1:0] out_474;
wire [32*C_WIDTH-1:0] out_475;
wire [32*C_WIDTH-1:0] out_476;
wire [32*C_WIDTH-1:0] out_477;
wire [32*C_WIDTH-1:0] out_478;
wire [32*C_WIDTH-1:0] out_479;
wire [32*C_WIDTH-1:0] out_480;
wire [32*C_WIDTH-1:0] out_481;
wire [32*C_WIDTH-1:0] out_482;
wire [32*C_WIDTH-1:0] out_483;
wire [32*C_WIDTH-1:0] out_484;
wire [32*C_WIDTH-1:0] out_485;
wire [32*C_WIDTH-1:0] out_486;
wire [32*C_WIDTH-1:0] out_487;
wire [32*C_WIDTH-1:0] out_488;
wire [32*C_WIDTH-1:0] out_489;
wire [32*C_WIDTH-1:0] out_490;
wire [32*C_WIDTH-1:0] out_491;
wire [32*C_WIDTH-1:0] out_492;
wire [32*C_WIDTH-1:0] out_493;
wire [32*C_WIDTH-1:0] out_494;
wire [32*C_WIDTH-1:0] out_495;
wire [32*C_WIDTH-1:0] out_496;
wire [32*C_WIDTH-1:0] out_497;
wire [32*C_WIDTH-1:0] out_498;
wire [32*C_WIDTH-1:0] out_499;
wire [32*C_WIDTH-1:0] out_500;
wire [32*C_WIDTH-1:0] out_501;
wire [32*C_WIDTH-1:0] out_502;
wire [32*C_WIDTH-1:0] out_503;
wire [32*C_WIDTH-1:0] out_504;
wire [32*C_WIDTH-1:0] out_505;
wire [32*C_WIDTH-1:0] out_506;
wire [32*C_WIDTH-1:0] out_507;
wire [32*C_WIDTH-1:0] out_508;
wire [32*C_WIDTH-1:0] out_509;
wire [32*C_WIDTH-1:0] out_510;
wire [32*C_WIDTH-1:0] out_511;
assign {act_0,act_1} = activation;
assign {weight_0,weight_1} = weight;

SA64 SA64_0 (.clk(clk),.rstn(rstn),.activation(act_0),.weight(weight_0),.out_act(act0_1),.out_weight(weight0_2),.control(control),
.c_out0(out_0),
.c_out1(out_1),
.c_out2(out_2),
.c_out3(out_3),
.c_out4(out_4),
.c_out5(out_5),
.c_out6(out_6),
.c_out7(out_7),
.c_out8(out_8),
.c_out9(out_9),
.c_out10(out_10),
.c_out11(out_11),
.c_out12(out_12),
.c_out13(out_13),
.c_out14(out_14),
.c_out15(out_15),
.c_out16(out_16),
.c_out17(out_17),
.c_out18(out_18),
.c_out19(out_19),
.c_out20(out_20),
.c_out21(out_21),
.c_out22(out_22),
.c_out23(out_23),
.c_out24(out_24),
.c_out25(out_25),
.c_out26(out_26),
.c_out27(out_27),
.c_out28(out_28),
.c_out29(out_29),
.c_out30(out_30),
.c_out31(out_31),
.c_out32(out_32),
.c_out33(out_33),
.c_out34(out_34),
.c_out35(out_35),
.c_out36(out_36),
.c_out37(out_37),
.c_out38(out_38),
.c_out39(out_39),
.c_out40(out_40),
.c_out41(out_41),
.c_out42(out_42),
.c_out43(out_43),
.c_out44(out_44),
.c_out45(out_45),
.c_out46(out_46),
.c_out47(out_47),
.c_out48(out_48),
.c_out49(out_49),
.c_out50(out_50),
.c_out51(out_51),
.c_out52(out_52),
.c_out53(out_53),
.c_out54(out_54),
.c_out55(out_55),
.c_out56(out_56),
.c_out57(out_57),
.c_out58(out_58),
.c_out59(out_59),
.c_out60(out_60),
.c_out61(out_61),
.c_out62(out_62),
.c_out63(out_63),
.c_out64(out_64),
.c_out65(out_65),
.c_out66(out_66),
.c_out67(out_67),
.c_out68(out_68),
.c_out69(out_69),
.c_out70(out_70),
.c_out71(out_71),
.c_out72(out_72),
.c_out73(out_73),
.c_out74(out_74),
.c_out75(out_75),
.c_out76(out_76),
.c_out77(out_77),
.c_out78(out_78),
.c_out79(out_79),
.c_out80(out_80),
.c_out81(out_81),
.c_out82(out_82),
.c_out83(out_83),
.c_out84(out_84),
.c_out85(out_85),
.c_out86(out_86),
.c_out87(out_87),
.c_out88(out_88),
.c_out89(out_89),
.c_out90(out_90),
.c_out91(out_91),
.c_out92(out_92),
.c_out93(out_93),
.c_out94(out_94),
.c_out95(out_95),
.c_out96(out_96),
.c_out97(out_97),
.c_out98(out_98),
.c_out99(out_99),
.c_out100(out_100),
.c_out101(out_101),
.c_out102(out_102),
.c_out103(out_103),
.c_out104(out_104),
.c_out105(out_105),
.c_out106(out_106),
.c_out107(out_107),
.c_out108(out_108),
.c_out109(out_109),
.c_out110(out_110),
.c_out111(out_111),
.c_out112(out_112),
.c_out113(out_113),
.c_out114(out_114),
.c_out115(out_115),
.c_out116(out_116),
.c_out117(out_117),
.c_out118(out_118),
.c_out119(out_119),
.c_out120(out_120),
.c_out121(out_121),
.c_out122(out_122),
.c_out123(out_123),
.c_out124(out_124),
.c_out125(out_125),
.c_out126(out_126),
.c_out127(out_127));
SA64 SA64_1 (.clk(clk),.rstn(rstn),.activation(act0_1),.weight(weight_1),.out_act(outact_0),.out_weight(weight1_3),.control(control),.c_out0(out_128),
.c_out1(out_129),
.c_out2(out_130),
.c_out3(out_131),
.c_out4(out_132),
.c_out5(out_133),
.c_out6(out_134),
.c_out7(out_135),
.c_out8(out_136),
.c_out9(out_137),
.c_out10(out_138),
.c_out11(out_139),
.c_out12(out_140),
.c_out13(out_141),
.c_out14(out_142),
.c_out15(out_143),
.c_out16(out_144),
.c_out17(out_145),
.c_out18(out_146),
.c_out19(out_147),
.c_out20(out_148),
.c_out21(out_149),
.c_out22(out_150),
.c_out23(out_151),
.c_out24(out_152),
.c_out25(out_153),
.c_out26(out_154),
.c_out27(out_155),
.c_out28(out_156),
.c_out29(out_157),
.c_out30(out_158),
.c_out31(out_159),
.c_out32(out_160),
.c_out33(out_161),
.c_out34(out_162),
.c_out35(out_163),
.c_out36(out_164),
.c_out37(out_165),
.c_out38(out_166),
.c_out39(out_167),
.c_out40(out_168),
.c_out41(out_169),
.c_out42(out_170),
.c_out43(out_171),
.c_out44(out_172),
.c_out45(out_173),
.c_out46(out_174),
.c_out47(out_175),
.c_out48(out_176),
.c_out49(out_177),
.c_out50(out_178),
.c_out51(out_179),
.c_out52(out_180),
.c_out53(out_181),
.c_out54(out_182),
.c_out55(out_183),
.c_out56(out_184),
.c_out57(out_185),
.c_out58(out_186),
.c_out59(out_187),
.c_out60(out_188),
.c_out61(out_189),
.c_out62(out_190),
.c_out63(out_191),
.c_out64(out_192),
.c_out65(out_193),
.c_out66(out_194),
.c_out67(out_195),
.c_out68(out_196),
.c_out69(out_197),
.c_out70(out_198),
.c_out71(out_199),
.c_out72(out_200),
.c_out73(out_201),
.c_out74(out_202),
.c_out75(out_203),
.c_out76(out_204),
.c_out77(out_205),
.c_out78(out_206),
.c_out79(out_207),
.c_out80(out_208),
.c_out81(out_209),
.c_out82(out_210),
.c_out83(out_211),
.c_out84(out_212),
.c_out85(out_213),
.c_out86(out_214),
.c_out87(out_215),
.c_out88(out_216),
.c_out89(out_217),
.c_out90(out_218),
.c_out91(out_219),
.c_out92(out_220),
.c_out93(out_221),
.c_out94(out_222),
.c_out95(out_223),
.c_out96(out_224),
.c_out97(out_225),
.c_out98(out_226),
.c_out99(out_227),
.c_out100(out_228),
.c_out101(out_229),
.c_out102(out_230),
.c_out103(out_231),
.c_out104(out_232),
.c_out105(out_233),
.c_out106(out_234),
.c_out107(out_235),
.c_out108(out_236),
.c_out109(out_237),
.c_out110(out_238),
.c_out111(out_239),
.c_out112(out_240),
.c_out113(out_241),
.c_out114(out_242),
.c_out115(out_243),
.c_out116(out_244),
.c_out117(out_245),
.c_out118(out_246),
.c_out119(out_247),
.c_out120(out_248),
.c_out121(out_249),
.c_out122(out_250),
.c_out123(out_251),
.c_out124(out_252),
.c_out125(out_253),
.c_out126(out_254),
.c_out127(out_255));
SA64 SA64_2 (.clk(clk),.rstn(rstn),.activation(act_1),.weight(weight0_2),.out_act(act2_3),.out_weight(outweight_0),.control(control),.c_out0(out_256),
.c_out1(out_257),
.c_out2(out_258),
.c_out3(out_259),
.c_out4(out_260),
.c_out5(out_261),
.c_out6(out_262),
.c_out7(out_263),
.c_out8(out_264),
.c_out9(out_265),
.c_out10(out_266),
.c_out11(out_267),
.c_out12(out_268),
.c_out13(out_269),
.c_out14(out_270),
.c_out15(out_271),
.c_out16(out_272),
.c_out17(out_273),
.c_out18(out_274),
.c_out19(out_275),
.c_out20(out_276),
.c_out21(out_277),
.c_out22(out_278),
.c_out23(out_279),
.c_out24(out_280),
.c_out25(out_281),
.c_out26(out_282),
.c_out27(out_283),
.c_out28(out_284),
.c_out29(out_285),
.c_out30(out_286),
.c_out31(out_287),
.c_out32(out_288),
.c_out33(out_289),
.c_out34(out_290),
.c_out35(out_291),
.c_out36(out_292),
.c_out37(out_293),
.c_out38(out_294),
.c_out39(out_295),
.c_out40(out_296),
.c_out41(out_297),
.c_out42(out_298),
.c_out43(out_299),
.c_out44(out_300),
.c_out45(out_301),
.c_out46(out_302),
.c_out47(out_303),
.c_out48(out_304),
.c_out49(out_305),
.c_out50(out_306),
.c_out51(out_307),
.c_out52(out_308),
.c_out53(out_309),
.c_out54(out_310),
.c_out55(out_311),
.c_out56(out_312),
.c_out57(out_313),
.c_out58(out_314),
.c_out59(out_315),
.c_out60(out_316),
.c_out61(out_317),
.c_out62(out_318),
.c_out63(out_319),
.c_out64(out_320),
.c_out65(out_321),
.c_out66(out_322),
.c_out67(out_323),
.c_out68(out_324),
.c_out69(out_325),
.c_out70(out_326),
.c_out71(out_327),
.c_out72(out_328),
.c_out73(out_329),
.c_out74(out_330),
.c_out75(out_331),
.c_out76(out_332),
.c_out77(out_333),
.c_out78(out_334),
.c_out79(out_335),
.c_out80(out_336),
.c_out81(out_337),
.c_out82(out_338),
.c_out83(out_339),
.c_out84(out_340),
.c_out85(out_341),
.c_out86(out_342),
.c_out87(out_343),
.c_out88(out_344),
.c_out89(out_345),
.c_out90(out_346),
.c_out91(out_347),
.c_out92(out_348),
.c_out93(out_349),
.c_out94(out_350),
.c_out95(out_351),
.c_out96(out_352),
.c_out97(out_353),
.c_out98(out_354),
.c_out99(out_355),
.c_out100(out_356),
.c_out101(out_357),
.c_out102(out_358),
.c_out103(out_359),
.c_out104(out_360),
.c_out105(out_361),
.c_out106(out_362),
.c_out107(out_363),
.c_out108(out_364),
.c_out109(out_365),
.c_out110(out_366),
.c_out111(out_367),
.c_out112(out_368),
.c_out113(out_369),
.c_out114(out_370),
.c_out115(out_371),
.c_out116(out_372),
.c_out117(out_373),
.c_out118(out_374),
.c_out119(out_375),
.c_out120(out_376),
.c_out121(out_377),
.c_out122(out_378),
.c_out123(out_379),
.c_out124(out_380),
.c_out125(out_381),
.c_out126(out_382),
.c_out127(out_383));
SA64 SA64_3 (.clk(clk),.rstn(rstn),.activation(act2_3),.weight(weight1_3),.out_act(outact_1),.out_weight(outweight_1),.control(control),.c_out0(out_384),
.c_out1(out_385),
.c_out2(out_386),
.c_out3(out_387),
.c_out4(out_388),
.c_out5(out_389),
.c_out6(out_390),
.c_out7(out_391),
.c_out8(out_392),
.c_out9(out_393),
.c_out10(out_394),
.c_out11(out_395),
.c_out12(out_396),
.c_out13(out_397),
.c_out14(out_398),
.c_out15(out_399),
.c_out16(out_400),
.c_out17(out_401),
.c_out18(out_402),
.c_out19(out_403),
.c_out20(out_404),
.c_out21(out_405),
.c_out22(out_406),
.c_out23(out_407),
.c_out24(out_408),
.c_out25(out_409),
.c_out26(out_410),
.c_out27(out_411),
.c_out28(out_412),
.c_out29(out_413),
.c_out30(out_414),
.c_out31(out_415),
.c_out32(out_416),
.c_out33(out_417),
.c_out34(out_418),
.c_out35(out_419),
.c_out36(out_420),
.c_out37(out_421),
.c_out38(out_422),
.c_out39(out_423),
.c_out40(out_424),
.c_out41(out_425),
.c_out42(out_426),
.c_out43(out_427),
.c_out44(out_428),
.c_out45(out_429),
.c_out46(out_430),
.c_out47(out_431),
.c_out48(out_432),
.c_out49(out_433),
.c_out50(out_434),
.c_out51(out_435),
.c_out52(out_436),
.c_out53(out_437),
.c_out54(out_438),
.c_out55(out_439),
.c_out56(out_440),
.c_out57(out_441),
.c_out58(out_442),
.c_out59(out_443),
.c_out60(out_444),
.c_out61(out_445),
.c_out62(out_446),
.c_out63(out_447),
.c_out64(out_448),
.c_out65(out_449),
.c_out66(out_450),
.c_out67(out_451),
.c_out68(out_452),
.c_out69(out_453),
.c_out70(out_454),
.c_out71(out_455),
.c_out72(out_456),
.c_out73(out_457),
.c_out74(out_458),
.c_out75(out_459),
.c_out76(out_460),
.c_out77(out_461),
.c_out78(out_462),
.c_out79(out_463),
.c_out80(out_464),
.c_out81(out_465),
.c_out82(out_466),
.c_out83(out_467),
.c_out84(out_468),
.c_out85(out_469),
.c_out86(out_470),
.c_out87(out_471),
.c_out88(out_472),
.c_out89(out_473),
.c_out90(out_474),
.c_out91(out_475),
.c_out92(out_476),
.c_out93(out_477),
.c_out94(out_478),
.c_out95(out_479),
.c_out96(out_480),
.c_out97(out_481),
.c_out98(out_482),
.c_out99(out_483),
.c_out100(out_484),
.c_out101(out_485),
.c_out102(out_486),
.c_out103(out_487),
.c_out104(out_488),
.c_out105(out_489),
.c_out106(out_490),
.c_out107(out_491),
.c_out108(out_492),
.c_out109(out_493),
.c_out110(out_494),
.c_out111(out_495),
.c_out112(out_496),
.c_out113(out_497),
.c_out114(out_498),
.c_out115(out_499),
.c_out116(out_500),
.c_out117(out_501),
.c_out118(out_502),
.c_out119(out_503),
.c_out120(out_504),
.c_out121(out_505),
.c_out122(out_506),
.c_out123(out_507),
.c_out124(out_508),
.c_out125(out_509),
.c_out126(out_510),
.c_out127(out_511));

assign out_act = {outact_0,outact_1};
assign out_weight = {outweight_0,outweight_1};

assign c_out0 = out_0;
assign c_out1 = out_1;
assign c_out2 = out_2;
assign c_out3 = out_3;
assign c_out4 = out_4;
assign c_out5 = out_5;
assign c_out6 = out_6;
assign c_out7 = out_7;
assign c_out8 = out_8;
assign c_out9 = out_9;
assign c_out10 = out_10;
assign c_out11 = out_11;
assign c_out12 = out_12;
assign c_out13 = out_13;
assign c_out14 = out_14;
assign c_out15 = out_15;
assign c_out16 = out_16;
assign c_out17 = out_17;
assign c_out18 = out_18;
assign c_out19 = out_19;
assign c_out20 = out_20;
assign c_out21 = out_21;
assign c_out22 = out_22;
assign c_out23 = out_23;
assign c_out24 = out_24;
assign c_out25 = out_25;
assign c_out26 = out_26;
assign c_out27 = out_27;
assign c_out28 = out_28;
assign c_out29 = out_29;
assign c_out30 = out_30;
assign c_out31 = out_31;
assign c_out32 = out_32;
assign c_out33 = out_33;
assign c_out34 = out_34;
assign c_out35 = out_35;
assign c_out36 = out_36;
assign c_out37 = out_37;
assign c_out38 = out_38;
assign c_out39 = out_39;
assign c_out40 = out_40;
assign c_out41 = out_41;
assign c_out42 = out_42;
assign c_out43 = out_43;
assign c_out44 = out_44;
assign c_out45 = out_45;
assign c_out46 = out_46;
assign c_out47 = out_47;
assign c_out48 = out_48;
assign c_out49 = out_49;
assign c_out50 = out_50;
assign c_out51 = out_51;
assign c_out52 = out_52;
assign c_out53 = out_53;
assign c_out54 = out_54;
assign c_out55 = out_55;
assign c_out56 = out_56;
assign c_out57 = out_57;
assign c_out58 = out_58;
assign c_out59 = out_59;
assign c_out60 = out_60;
assign c_out61 = out_61;
assign c_out62 = out_62;
assign c_out63 = out_63;
assign c_out64 = out_64;
assign c_out65 = out_65;
assign c_out66 = out_66;
assign c_out67 = out_67;
assign c_out68 = out_68;
assign c_out69 = out_69;
assign c_out70 = out_70;
assign c_out71 = out_71;
assign c_out72 = out_72;
assign c_out73 = out_73;
assign c_out74 = out_74;
assign c_out75 = out_75;
assign c_out76 = out_76;
assign c_out77 = out_77;
assign c_out78 = out_78;
assign c_out79 = out_79;
assign c_out80 = out_80;
assign c_out81 = out_81;
assign c_out82 = out_82;
assign c_out83 = out_83;
assign c_out84 = out_84;
assign c_out85 = out_85;
assign c_out86 = out_86;
assign c_out87 = out_87;
assign c_out88 = out_88;
assign c_out89 = out_89;
assign c_out90 = out_90;
assign c_out91 = out_91;
assign c_out92 = out_92;
assign c_out93 = out_93;
assign c_out94 = out_94;
assign c_out95 = out_95;
assign c_out96 = out_96;
assign c_out97 = out_97;
assign c_out98 = out_98;
assign c_out99 = out_99;
assign c_out100 = out_100;
assign c_out101 = out_101;
assign c_out102 = out_102;
assign c_out103 = out_103;
assign c_out104 = out_104;
assign c_out105 = out_105;
assign c_out106 = out_106;
assign c_out107 = out_107;
assign c_out108 = out_108;
assign c_out109 = out_109;
assign c_out110 = out_110;
assign c_out111 = out_111;
assign c_out112 = out_112;
assign c_out113 = out_113;
assign c_out114 = out_114;
assign c_out115 = out_115;
assign c_out116 = out_116;
assign c_out117 = out_117;
assign c_out118 = out_118;
assign c_out119 = out_119;
assign c_out120 = out_120;
assign c_out121 = out_121;
assign c_out122 = out_122;
assign c_out123 = out_123;
assign c_out124 = out_124;
assign c_out125 = out_125;
assign c_out126 = out_126;
assign c_out127 = out_127;
assign c_out128 = out_128;
assign c_out129 = out_129;
assign c_out130 = out_130;
assign c_out131 = out_131;
assign c_out132 = out_132;
assign c_out133 = out_133;
assign c_out134 = out_134;
assign c_out135 = out_135;
assign c_out136 = out_136;
assign c_out137 = out_137;
assign c_out138 = out_138;
assign c_out139 = out_139;
assign c_out140 = out_140;
assign c_out141 = out_141;
assign c_out142 = out_142;
assign c_out143 = out_143;
assign c_out144 = out_144;
assign c_out145 = out_145;
assign c_out146 = out_146;
assign c_out147 = out_147;
assign c_out148 = out_148;
assign c_out149 = out_149;
assign c_out150 = out_150;
assign c_out151 = out_151;
assign c_out152 = out_152;
assign c_out153 = out_153;
assign c_out154 = out_154;
assign c_out155 = out_155;
assign c_out156 = out_156;
assign c_out157 = out_157;
assign c_out158 = out_158;
assign c_out159 = out_159;
assign c_out160 = out_160;
assign c_out161 = out_161;
assign c_out162 = out_162;
assign c_out163 = out_163;
assign c_out164 = out_164;
assign c_out165 = out_165;
assign c_out166 = out_166;
assign c_out167 = out_167;
assign c_out168 = out_168;
assign c_out169 = out_169;
assign c_out170 = out_170;
assign c_out171 = out_171;
assign c_out172 = out_172;
assign c_out173 = out_173;
assign c_out174 = out_174;
assign c_out175 = out_175;
assign c_out176 = out_176;
assign c_out177 = out_177;
assign c_out178 = out_178;
assign c_out179 = out_179;
assign c_out180 = out_180;
assign c_out181 = out_181;
assign c_out182 = out_182;
assign c_out183 = out_183;
assign c_out184 = out_184;
assign c_out185 = out_185;
assign c_out186 = out_186;
assign c_out187 = out_187;
assign c_out188 = out_188;
assign c_out189 = out_189;
assign c_out190 = out_190;
assign c_out191 = out_191;
assign c_out192 = out_192;
assign c_out193 = out_193;
assign c_out194 = out_194;
assign c_out195 = out_195;
assign c_out196 = out_196;
assign c_out197 = out_197;
assign c_out198 = out_198;
assign c_out199 = out_199;
assign c_out200 = out_200;
assign c_out201 = out_201;
assign c_out202 = out_202;
assign c_out203 = out_203;
assign c_out204 = out_204;
assign c_out205 = out_205;
assign c_out206 = out_206;
assign c_out207 = out_207;
assign c_out208 = out_208;
assign c_out209 = out_209;
assign c_out210 = out_210;
assign c_out211 = out_211;
assign c_out212 = out_212;
assign c_out213 = out_213;
assign c_out214 = out_214;
assign c_out215 = out_215;
assign c_out216 = out_216;
assign c_out217 = out_217;
assign c_out218 = out_218;
assign c_out219 = out_219;
assign c_out220 = out_220;
assign c_out221 = out_221;
assign c_out222 = out_222;
assign c_out223 = out_223;
assign c_out224 = out_224;
assign c_out225 = out_225;
assign c_out226 = out_226;
assign c_out227 = out_227;
assign c_out228 = out_228;
assign c_out229 = out_229;
assign c_out230 = out_230;
assign c_out231 = out_231;
assign c_out232 = out_232;
assign c_out233 = out_233;
assign c_out234 = out_234;
assign c_out235 = out_235;
assign c_out236 = out_236;
assign c_out237 = out_237;
assign c_out238 = out_238;
assign c_out239 = out_239;
assign c_out240 = out_240;
assign c_out241 = out_241;
assign c_out242 = out_242;
assign c_out243 = out_243;
assign c_out244 = out_244;
assign c_out245 = out_245;
assign c_out246 = out_246;
assign c_out247 = out_247;
assign c_out248 = out_248;
assign c_out249 = out_249;
assign c_out250 = out_250;
assign c_out251 = out_251;
assign c_out252 = out_252;
assign c_out253 = out_253;
assign c_out254 = out_254;
assign c_out255 = out_255;
assign c_out256 = out_256;
assign c_out257 = out_257;
assign c_out258 = out_258;
assign c_out259 = out_259;
assign c_out260 = out_260;
assign c_out261 = out_261;
assign c_out262 = out_262;
assign c_out263 = out_263;
assign c_out264 = out_264;
assign c_out265 = out_265;
assign c_out266 = out_266;
assign c_out267 = out_267;
assign c_out268 = out_268;
assign c_out269 = out_269;
assign c_out270 = out_270;
assign c_out271 = out_271;
assign c_out272 = out_272;
assign c_out273 = out_273;
assign c_out274 = out_274;
assign c_out275 = out_275;
assign c_out276 = out_276;
assign c_out277 = out_277;
assign c_out278 = out_278;
assign c_out279 = out_279;
assign c_out280 = out_280;
assign c_out281 = out_281;
assign c_out282 = out_282;
assign c_out283 = out_283;
assign c_out284 = out_284;
assign c_out285 = out_285;
assign c_out286 = out_286;
assign c_out287 = out_287;
assign c_out288 = out_288;
assign c_out289 = out_289;
assign c_out290 = out_290;
assign c_out291 = out_291;
assign c_out292 = out_292;
assign c_out293 = out_293;
assign c_out294 = out_294;
assign c_out295 = out_295;
assign c_out296 = out_296;
assign c_out297 = out_297;
assign c_out298 = out_298;
assign c_out299 = out_299;
assign c_out300 = out_300;
assign c_out301 = out_301;
assign c_out302 = out_302;
assign c_out303 = out_303;
assign c_out304 = out_304;
assign c_out305 = out_305;
assign c_out306 = out_306;
assign c_out307 = out_307;
assign c_out308 = out_308;
assign c_out309 = out_309;
assign c_out310 = out_310;
assign c_out311 = out_311;
assign c_out312 = out_312;
assign c_out313 = out_313;
assign c_out314 = out_314;
assign c_out315 = out_315;
assign c_out316 = out_316;
assign c_out317 = out_317;
assign c_out318 = out_318;
assign c_out319 = out_319;
assign c_out320 = out_320;
assign c_out321 = out_321;
assign c_out322 = out_322;
assign c_out323 = out_323;
assign c_out324 = out_324;
assign c_out325 = out_325;
assign c_out326 = out_326;
assign c_out327 = out_327;
assign c_out328 = out_328;
assign c_out329 = out_329;
assign c_out330 = out_330;
assign c_out331 = out_331;
assign c_out332 = out_332;
assign c_out333 = out_333;
assign c_out334 = out_334;
assign c_out335 = out_335;
assign c_out336 = out_336;
assign c_out337 = out_337;
assign c_out338 = out_338;
assign c_out339 = out_339;
assign c_out340 = out_340;
assign c_out341 = out_341;
assign c_out342 = out_342;
assign c_out343 = out_343;
assign c_out344 = out_344;
assign c_out345 = out_345;
assign c_out346 = out_346;
assign c_out347 = out_347;
assign c_out348 = out_348;
assign c_out349 = out_349;
assign c_out350 = out_350;
assign c_out351 = out_351;
assign c_out352 = out_352;
assign c_out353 = out_353;
assign c_out354 = out_354;
assign c_out355 = out_355;
assign c_out356 = out_356;
assign c_out357 = out_357;
assign c_out358 = out_358;
assign c_out359 = out_359;
assign c_out360 = out_360;
assign c_out361 = out_361;
assign c_out362 = out_362;
assign c_out363 = out_363;
assign c_out364 = out_364;
assign c_out365 = out_365;
assign c_out366 = out_366;
assign c_out367 = out_367;
assign c_out368 = out_368;
assign c_out369 = out_369;
assign c_out370 = out_370;
assign c_out371 = out_371;
assign c_out372 = out_372;
assign c_out373 = out_373;
assign c_out374 = out_374;
assign c_out375 = out_375;
assign c_out376 = out_376;
assign c_out377 = out_377;
assign c_out378 = out_378;
assign c_out379 = out_379;
assign c_out380 = out_380;
assign c_out381 = out_381;
assign c_out382 = out_382;
assign c_out383 = out_383;
assign c_out384 = out_384;
assign c_out385 = out_385;
assign c_out386 = out_386;
assign c_out387 = out_387;
assign c_out388 = out_388;
assign c_out389 = out_389;
assign c_out390 = out_390;
assign c_out391 = out_391;
assign c_out392 = out_392;
assign c_out393 = out_393;
assign c_out394 = out_394;
assign c_out395 = out_395;
assign c_out396 = out_396;
assign c_out397 = out_397;
assign c_out398 = out_398;
assign c_out399 = out_399;
assign c_out400 = out_400;
assign c_out401 = out_401;
assign c_out402 = out_402;
assign c_out403 = out_403;
assign c_out404 = out_404;
assign c_out405 = out_405;
assign c_out406 = out_406;
assign c_out407 = out_407;
assign c_out408 = out_408;
assign c_out409 = out_409;
assign c_out410 = out_410;
assign c_out411 = out_411;
assign c_out412 = out_412;
assign c_out413 = out_413;
assign c_out414 = out_414;
assign c_out415 = out_415;
assign c_out416 = out_416;
assign c_out417 = out_417;
assign c_out418 = out_418;
assign c_out419 = out_419;
assign c_out420 = out_420;
assign c_out421 = out_421;
assign c_out422 = out_422;
assign c_out423 = out_423;
assign c_out424 = out_424;
assign c_out425 = out_425;
assign c_out426 = out_426;
assign c_out427 = out_427;
assign c_out428 = out_428;
assign c_out429 = out_429;
assign c_out430 = out_430;
assign c_out431 = out_431;
assign c_out432 = out_432;
assign c_out433 = out_433;
assign c_out434 = out_434;
assign c_out435 = out_435;
assign c_out436 = out_436;
assign c_out437 = out_437;
assign c_out438 = out_438;
assign c_out439 = out_439;
assign c_out440 = out_440;
assign c_out441 = out_441;
assign c_out442 = out_442;
assign c_out443 = out_443;
assign c_out444 = out_444;
assign c_out445 = out_445;
assign c_out446 = out_446;
assign c_out447 = out_447;
assign c_out448 = out_448;
assign c_out449 = out_449;
assign c_out450 = out_450;
assign c_out451 = out_451;
assign c_out452 = out_452;
assign c_out453 = out_453;
assign c_out454 = out_454;
assign c_out455 = out_455;
assign c_out456 = out_456;
assign c_out457 = out_457;
assign c_out458 = out_458;
assign c_out459 = out_459;
assign c_out460 = out_460;
assign c_out461 = out_461;
assign c_out462 = out_462;
assign c_out463 = out_463;
assign c_out464 = out_464;
assign c_out465 = out_465;
assign c_out466 = out_466;
assign c_out467 = out_467;
assign c_out468 = out_468;
assign c_out469 = out_469;
assign c_out470 = out_470;
assign c_out471 = out_471;
assign c_out472 = out_472;
assign c_out473 = out_473;
assign c_out474 = out_474;
assign c_out475 = out_475;
assign c_out476 = out_476;
assign c_out477 = out_477;
assign c_out478 = out_478;
assign c_out479 = out_479;
assign c_out480 = out_480;
assign c_out481 = out_481;
assign c_out482 = out_482;
assign c_out483 = out_483;
assign c_out484 = out_484;
assign c_out485 = out_485;
assign c_out486 = out_486;
assign c_out487 = out_487;
assign c_out488 = out_488;
assign c_out489 = out_489;
assign c_out490 = out_490;
assign c_out491 = out_491;
assign c_out492 = out_492;
assign c_out493 = out_493;
assign c_out494 = out_494;
assign c_out495 = out_495;
assign c_out496 = out_496;
assign c_out497 = out_497;
assign c_out498 = out_498;
assign c_out499 = out_499;
assign c_out500 = out_500;
assign c_out501 = out_501;
assign c_out502 = out_502;
assign c_out503 = out_503;
assign c_out504 = out_504;
assign c_out505 = out_505;
assign c_out506 = out_506;
assign c_out507 = out_507;
assign c_out508 = out_508;
assign c_out509 = out_509;
assign c_out510 = out_510;
assign c_out511 = out_511;
​


endmodule
